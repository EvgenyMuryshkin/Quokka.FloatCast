/*
 *  Float to 64 bit integer converter
 *
 *  Copyright (C) 2019  Evgeny Muryshkin <evmuryshkin@gmail.com>
 *
 *  Part of Quokka FPGA toolkit
 *  https://github.com/EvgenyMuryshkin/QuokkaEvaluation
 *
 *  Permission to use, copy, modify, and/or distribute this software for any
 *  purpose with or without fee is hereby granted, provided that the above
 *  copyright notice and this permission notice appear in all copies.
 *
 *  THE SOFTWARE IS PROVIDED "AS IS" AND THE AUTHOR DISCLAIMS ALL WARRANTIES
 *  WITH REGARD TO THIS SOFTWARE INCLUDING ALL IMPLIED WARRANTIES OF
 *  MERCHANTABILITY AND FITNESS. IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR
 *  ANY SPECIAL, DIRECT, INDIRECT, OR CONSEQUENTIAL DAMAGES OR ANY DAMAGES
 *  WHATSOEVER RESULTING FROM LOSS OF USE, DATA OR PROFITS, WHETHER IN AN
 *  ACTION OF CONTRACT, NEGLIGENCE OR OTHER TORTIOUS ACTION, ARISING OUT OF
 *  OR IN CONNECTION WITH THE USE OR PERFORMANCE OF THIS SOFTWARE.
 */
import uvm_pkg::*;
`include "uvm_macros.svh"

//---------------------------------------
// Interface for the FloatToInt DUT
//---------------------------------------
interface FloatToInt_IF(
	input bit clk,
  	input inTrigger,
  	input [31:0] inData,
  	input [63:0] outData,
	input outReady,
  	input outException
);

  clocking cb @(posedge clk);
    output     inTrigger;
    output     inData;
    input    outData;
    input    outReady;
    input    outException;
  endclocking // cb

endinterface: FloatToInt_IF

//---------------
// Interface bind
//---------------
bind FloatToInt FloatToInt_IF FloatToInt_IF0(
  .clk(clk),
  .inTrigger(inTrigger),
  .inData(inData),
  .outData(outData),
  .outReady(outReady),
  .outException(outException)
);

//----------------
// environment env
//----------------
class env extends uvm_env;

  virtual FloatToInt_IF m_if;

  function new(string name, uvm_component parent = null);
    super.new(name, parent);
  endfunction
  
  function void connect_phase(uvm_phase phase);
    `uvm_info("LABEL", "Started connect phase.", UVM_HIGH);
    // Get the interface from the resource database.
    assert(uvm_resource_db#(virtual FloatToInt_IF)::read_by_name(
      get_full_name(), "FloatToInt_IF", m_if));
    `uvm_info("LABEL", "Finished connect phase.", UVM_HIGH);
  endfunction: connect_phase

  task fullCycle();
    begin
      repeat(2) @(m_if.cb);
    end
  endtask
  
  task convertSigned(int unsigned value, longint expected, string hint);
    begin
      m_if.cb.inData <= value;
      m_if.cb.inTrigger <= 1;
      fullCycle();
      
      m_if.cb.inTrigger <= 0;
      repeat(64) fullCycle();

      `uvm_info("RESULT", $sformatf("[Float Hex] %0x [Float Value] %s [Expecting] %0d [Actual] %0x", value, hint, expected, m_if.cb.outData), UVM_LOW);
      if (m_if.cb.outReady != 1)
        `uvm_error("outReady", "Did not finish convertion");
      
      if (m_if.cb.outData != expected)
        `uvm_error("outData", "Result did not match");

    end
  endtask
  
  task run_phase(uvm_phase phase);
    phase.raise_objection(this);
    `uvm_info("LABEL", "Started run phase.", UVM_HIGH);
    begin
      @(m_if.cb);
     
      convertSigned(32'hFFC00000, 64'h8000000000000000, "NaN"); // NaN
      convertSigned(32'hFF800000, 64'h8000000000000000, "Neg Inf"); // Neg Inf
      convertSigned(32'hDE800002, 64'hBFFFFF0000000000, "-4611687000000000000.000000"); // -4611687000000000000.000000
      convertSigned(32'hDE800001, 64'hBFFFFF8000000000, "-4611687000000000000.000000"); // -4611687000000000000.000000
      convertSigned(32'hDE800000, 64'hC000000000000000, "-4611686000000000000.000000"); // -4611686000000000000.000000
      convertSigned(32'hDE000002, 64'hDFFFFF8000000000, "-2305844000000000000.000000"); // -2305844000000000000.000000
      convertSigned(32'hDE000001, 64'hDFFFFFC000000000, "-2305843000000000000.000000"); // -2305843000000000000.000000
      convertSigned(32'hDE000000, 64'hE000000000000000, "-2305843000000000000.000000"); // -2305843000000000000.000000
      convertSigned(32'hDD800002, 64'hEFFFFFC000000000, "-1152922000000000000.000000"); // -1152922000000000000.000000
      convertSigned(32'hDD800001, 64'hEFFFFFE000000000, "-1152922000000000000.000000"); // -1152922000000000000.000000
      convertSigned(32'hDD800000, 64'hF000000000000000, "-1152922000000000000.000000"); // -1152922000000000000.000000
      convertSigned(32'hDD000002, 64'hF7FFFFE000000000, "-576460900000000000.000000"); // -576460900000000000.000000
      convertSigned(32'hDD000001, 64'hF7FFFFF000000000, "-576460800000000000.000000"); // -576460800000000000.000000
      convertSigned(32'hDD000000, 64'hF800000000000000, "-576460800000000000.000000"); // -576460800000000000.000000
      convertSigned(32'hDC800002, 64'hFBFFFFF000000000, "-288230400000000000.000000"); // -288230400000000000.000000
      convertSigned(32'hDC800001, 64'hFBFFFFF800000000, "-288230400000000000.000000"); // -288230400000000000.000000
      convertSigned(32'hDC800000, 64'hFC00000000000000, "-288230400000000000.000000"); // -288230400000000000.000000
      convertSigned(32'hDC000002, 64'hFDFFFFF800000000, "-144115200000000000.000000"); // -144115200000000000.000000
      convertSigned(32'hDC000001, 64'hFDFFFFFC00000000, "-144115200000000000.000000"); // -144115200000000000.000000
      convertSigned(32'hDC000000, 64'hFE00000000000000, "-144115200000000000.000000"); // -144115200000000000.000000
      convertSigned(32'hDB800002, 64'hFEFFFFFC00000000, "-72057610000000000.000000"); // -72057610000000000.000000
      convertSigned(32'hDB800001, 64'hFEFFFFFE00000000, "-72057600000000000.000000"); // -72057600000000000.000000
      convertSigned(32'hDB800000, 64'hFF00000000000000, "-72057590000000000.000000"); // -72057590000000000.000000
      convertSigned(32'hDB000002, 64'hFF7FFFFE00000000, "-36028810000000000.000000"); // -36028810000000000.000000
      convertSigned(32'hDB000001, 64'hFF7FFFFF00000000, "-36028800000000000.000000"); // -36028800000000000.000000
      convertSigned(32'hDB000000, 64'hFF80000000000000, "-36028800000000000.000000"); // -36028800000000000.000000
      convertSigned(32'hDA800002, 64'hFFBFFFFF00000000, "-18014400000000000.000000"); // -18014400000000000.000000
      convertSigned(32'hDA800001, 64'hFFBFFFFF80000000, "-18014400000000000.000000"); // -18014400000000000.000000
      convertSigned(32'hDA800000, 64'hFFC0000000000000, "-18014400000000000.000000"); // -18014400000000000.000000
      convertSigned(32'hDA000002, 64'hFFDFFFFF80000000, "-9007201000000000.000000"); // -9007201000000000.000000
      convertSigned(32'hDA000001, 64'hFFDFFFFFC0000000, "-9007200000000000.000000"); // -9007200000000000.000000
      convertSigned(32'hDA000000, 64'hFFE0000000000000, "-9007199000000000.000000"); // -9007199000000000.000000
      convertSigned(32'hD9800002, 64'hFFEFFFFFC0000000, "-4503601000000000.000000"); // -4503601000000000.000000
      convertSigned(32'hD9800001, 64'hFFEFFFFFE0000000, "-4503600000000000.000000"); // -4503600000000000.000000
      convertSigned(32'hD9800000, 64'hFFF0000000000000, "-4503600000000000.000000"); // -4503600000000000.000000
      convertSigned(32'hD9000002, 64'hFFF7FFFFE0000000, "-2251800000000000.000000"); // -2251800000000000.000000
      convertSigned(32'hD9000001, 64'hFFF7FFFFF0000000, "-2251800000000000.000000"); // -2251800000000000.000000
      convertSigned(32'hD9000000, 64'hFFF8000000000000, "-2251800000000000.000000"); // -2251800000000000.000000
      convertSigned(32'hD8800002, 64'hFFFBFFFFF0000000, "-1125900000000000.000000"); // -1125900000000000.000000
      convertSigned(32'hD8800001, 64'hFFFBFFFFF8000000, "-1125900000000000.000000"); // -1125900000000000.000000
      convertSigned(32'hD8800000, 64'hFFFC000000000000, "-1125900000000000.000000"); // -1125900000000000.000000
      convertSigned(32'hD8000002, 64'hFFFDFFFFF8000000, "-562950100000000.000000"); // -562950100000000.000000
      convertSigned(32'hD8000001, 64'hFFFDFFFFFC000000, "-562950000000000.000000"); // -562950000000000.000000
      convertSigned(32'hD8000000, 64'hFFFE000000000000, "-562950000000000.000000"); // -562950000000000.000000
      convertSigned(32'hD7800002, 64'hFFFEFFFFFC000000, "-281475000000000.000000"); // -281475000000000.000000
      convertSigned(32'hD7800001, 64'hFFFEFFFFFE000000, "-281475000000000.000000"); // -281475000000000.000000
      convertSigned(32'hD7800000, 64'hFFFF000000000000, "-281475000000000.000000"); // -281475000000000.000000
      convertSigned(32'hD7000002, 64'hFFFF7FFFFE000000, "-140737500000000.000000"); // -140737500000000.000000
      convertSigned(32'hD7000001, 64'hFFFF7FFFFF000000, "-140737500000000.000000"); // -140737500000000.000000
      convertSigned(32'hD7000000, 64'hFFFF800000000000, "-140737500000000.000000"); // -140737500000000.000000
      convertSigned(32'hD6800002, 64'hFFFFBFFFFF000000, "-70368760000000.000000"); // -70368760000000.000000
      convertSigned(32'hD6800001, 64'hFFFFBFFFFF800000, "-70368750000000.000000"); // -70368750000000.000000
      convertSigned(32'hD6800000, 64'hFFFFC00000000000, "-70368740000000.000000"); // -70368740000000.000000
      convertSigned(32'hD6000002, 64'hFFFFDFFFFF800000, "-35184380000000.000000"); // -35184380000000.000000
      convertSigned(32'hD6000001, 64'hFFFFDFFFFFC00000, "-35184380000000.000000"); // -35184380000000.000000
      convertSigned(32'hD6000000, 64'hFFFFE00000000000, "-35184370000000.000000"); // -35184370000000.000000
      convertSigned(32'hD5800002, 64'hFFFFEFFFFFC00000, "-17592190000000.000000"); // -17592190000000.000000
      convertSigned(32'hD5800001, 64'hFFFFEFFFFFE00000, "-17592190000000.000000"); // -17592190000000.000000
      convertSigned(32'hD5800000, 64'hFFFFF00000000000, "-17592190000000.000000"); // -17592190000000.000000
      convertSigned(32'hD5000002, 64'hFFFFF7FFFFE00000, "-8796095000000.000000"); // -8796095000000.000000
      convertSigned(32'hD5000001, 64'hFFFFF7FFFFF00000, "-8796094000000.000000"); // -8796094000000.000000
      convertSigned(32'hD5000000, 64'hFFFFF80000000000, "-8796093000000.000000"); // -8796093000000.000000
      convertSigned(32'hD4800002, 64'hFFFFFBFFFFF00000, "-4398048000000.000000"); // -4398048000000.000000
      convertSigned(32'hD4800001, 64'hFFFFFBFFFFF80000, "-4398047000000.000000"); // -4398047000000.000000
      convertSigned(32'hD4800000, 64'hFFFFFC0000000000, "-4398047000000.000000"); // -4398047000000.000000
      convertSigned(32'hD4000002, 64'hFFFFFDFFFFF80000, "-2199024000000.000000"); // -2199024000000.000000
      convertSigned(32'hD4000001, 64'hFFFFFDFFFFFC0000, "-2199024000000.000000"); // -2199024000000.000000
      convertSigned(32'hD4000000, 64'hFFFFFE0000000000, "-2199023000000.000000"); // -2199023000000.000000
      convertSigned(32'hD3800002, 64'hFFFFFEFFFFFC0000, "-1099512000000.000000"); // -1099512000000.000000
      convertSigned(32'hD3800001, 64'hFFFFFEFFFFFE0000, "-1099512000000.000000"); // -1099512000000.000000
      convertSigned(32'hD3800000, 64'hFFFFFF0000000000, "-1099512000000.000000"); // -1099512000000.000000
      convertSigned(32'hD3000002, 64'hFFFFFF7FFFFE0000, "-549755900000.000000"); // -549755900000.000000
      convertSigned(32'hD3000001, 64'hFFFFFF7FFFFF0000, "-549755900000.000000"); // -549755900000.000000
      convertSigned(32'hD3000000, 64'hFFFFFF8000000000, "-549755800000.000000"); // -549755800000.000000
      convertSigned(32'hD2800002, 64'hFFFFFFBFFFFF0000, "-274878000000.000000"); // -274878000000.000000
      convertSigned(32'hD2800001, 64'hFFFFFFBFFFFF8000, "-274877900000.000000"); // -274877900000.000000
      convertSigned(32'hD2800000, 64'hFFFFFFC000000000, "-274877900000.000000"); // -274877900000.000000
      convertSigned(32'hD2000002, 64'hFFFFFFDFFFFF8000, "-137439000000.000000"); // -137439000000.000000
      convertSigned(32'hD2000001, 64'hFFFFFFDFFFFFC000, "-137439000000.000000"); // -137439000000.000000
      convertSigned(32'hD2000000, 64'hFFFFFFE000000000, "-137439000000.000000"); // -137439000000.000000
      convertSigned(32'hD1800002, 64'hFFFFFFEFFFFFC000, "-68719490000.000000"); // -68719490000.000000
      convertSigned(32'hD1800001, 64'hFFFFFFEFFFFFE000, "-68719480000.000000"); // -68719480000.000000
      convertSigned(32'hD1800000, 64'hFFFFFFF000000000, "-68719480000.000000"); // -68719480000.000000
      convertSigned(32'hD1000002, 64'hFFFFFFF7FFFFE000, "-34359750000.000000"); // -34359750000.000000
      convertSigned(32'hD1000001, 64'hFFFFFFF7FFFFF000, "-34359740000.000000"); // -34359740000.000000
      convertSigned(32'hD1000000, 64'hFFFFFFF800000000, "-34359740000.000000"); // -34359740000.000000
      convertSigned(32'hD0800002, 64'hFFFFFFFBFFFFF000, "-17179870000.000000"); // -17179870000.000000
      convertSigned(32'hD0800001, 64'hFFFFFFFBFFFFF800, "-17179870000.000000"); // -17179870000.000000
      convertSigned(32'hD0800000, 64'hFFFFFFFC00000000, "-17179870000.000000"); // -17179870000.000000
      convertSigned(32'hD0000002, 64'hFFFFFFFDFFFFF800, "-8589937000.000000"); // -8589937000.000000
      convertSigned(32'hD0000001, 64'hFFFFFFFDFFFFFC00, "-8589936000.000000"); // -8589936000.000000
      convertSigned(32'hD0000000, 64'hFFFFFFFE00000000, "-8589935000.000000"); // -8589935000.000000
      convertSigned(32'hCF800002, 64'hFFFFFFFEFFFFFC00, "-4294968000.000000"); // -4294968000.000000
      convertSigned(32'hCF800001, 64'hFFFFFFFEFFFFFE00, "-4294968000.000000"); // -4294968000.000000
      convertSigned(32'hCF800000, 64'hFFFFFFFF00000000, "-4294967000.000000"); // -4294967000.000000
      convertSigned(32'hCF000002, 64'hFFFFFFFF7FFFFE00, "-2147484000.000000"); // -2147484000.000000
      convertSigned(32'hCF000001, 64'hFFFFFFFF7FFFFF00, "-2147484000.000000"); // -2147484000.000000
      convertSigned(32'hCF000000, 64'hFFFFFFFF80000000, "-2147484000.000000"); // -2147484000.000000
      convertSigned(32'hCE800002, 64'hFFFFFFFFBFFFFF00, "-1073742000.000000"); // -1073742000.000000
      convertSigned(32'hCE800001, 64'hFFFFFFFFBFFFFF80, "-1073742000.000000"); // -1073742000.000000
      convertSigned(32'hCE800000, 64'hFFFFFFFFC0000000, "-1073742000.000000"); // -1073742000.000000
      convertSigned(32'hCE000002, 64'hFFFFFFFFDFFFFF80, "-536871000.000000"); // -536871000.000000
      convertSigned(32'hCE000001, 64'hFFFFFFFFDFFFFFC0, "-536871000.000000"); // -536871000.000000
      convertSigned(32'hCE000000, 64'hFFFFFFFFE0000000, "-536870900.000000"); // -536870900.000000
      convertSigned(32'hCD800002, 64'hFFFFFFFFEFFFFFC0, "-268435500.000000"); // -268435500.000000
      convertSigned(32'hCD800001, 64'hFFFFFFFFEFFFFFE0, "-268435500.000000"); // -268435500.000000
      convertSigned(32'hCD800000, 64'hFFFFFFFFF0000000, "-268435500.000000"); // -268435500.000000
      convertSigned(32'hCD000002, 64'hFFFFFFFFF7FFFFE0, "-134217800.000000"); // -134217800.000000
      convertSigned(32'hCD000001, 64'hFFFFFFFFF7FFFFF0, "-134217700.000000"); // -134217700.000000
      convertSigned(32'hCD000000, 64'hFFFFFFFFF8000000, "-134217700.000000"); // -134217700.000000
      convertSigned(32'hCC800002, 64'hFFFFFFFFFBFFFFF0, "-67108880.000000"); // -67108880.000000
      convertSigned(32'hCC800001, 64'hFFFFFFFFFBFFFFF8, "-67108870.000000"); // -67108870.000000
      convertSigned(32'hCC800000, 64'hFFFFFFFFFC000000, "-67108860.000000"); // -67108860.000000
      convertSigned(32'hCC000002, 64'hFFFFFFFFFDFFFFF8, "-33554440.000000"); // -33554440.000000
      convertSigned(32'hCC000001, 64'hFFFFFFFFFDFFFFFC, "-33554440.000000"); // -33554440.000000
      convertSigned(32'hCC000000, 64'hFFFFFFFFFE000000, "-33554430.000000"); // -33554430.000000
      convertSigned(32'hCB800002, 64'hFFFFFFFFFEFFFFFC, "-16777220.000000"); // -16777220.000000
      convertSigned(32'hCB800001, 64'hFFFFFFFFFEFFFFFE, "-16777220.000000"); // -16777220.000000
      convertSigned(32'hCB800000, 64'hFFFFFFFFFF000000, "-16777220.000000"); // -16777220.000000
      convertSigned(32'hCB000001, 64'hFFFFFFFFFF7FFFFF, "-8388609"); // -8388609
      convertSigned(32'hCB000000, 64'hFFFFFFFFFF800000, "-8388608.000000"); // -8388608.000000
      convertSigned(32'hCAFFFFFF, 64'hFFFFFFFFFF800001, "-8388608.000000"); // -8388608.000000
      convertSigned(32'hCAFFFFFE, 64'hFFFFFFFFFF800001, "-8388607"); // -8388607
      convertSigned(32'hCAFFFFFD, 64'hFFFFFFFFFF800002, "-8388606.000000"); // -8388606.000000
      convertSigned(32'hCA800002, 64'hFFFFFFFFFFBFFFFF, "-4194305"); // -4194305
      convertSigned(32'hCA800001, 64'hFFFFFFFFFFC00000, "-4194304.000000"); // -4194304.000000
      convertSigned(32'hCA800000, 64'hFFFFFFFFFFC00000, "-4194304"); // -4194304
      convertSigned(32'hCA7FFFFE, 64'hFFFFFFFFFFC00001, "-4194304.000000"); // -4194304.000000
      convertSigned(32'hCA7FFFFC, 64'hFFFFFFFFFFC00001, "-4194303"); // -4194303
      convertSigned(32'hCA7FFFFA, 64'hFFFFFFFFFFC00002, "-4194302.000000"); // -4194302.000000
      convertSigned(32'hCA000004, 64'hFFFFFFFFFFDFFFFF, "-2097153"); // -2097153
      convertSigned(32'hCA000002, 64'hFFFFFFFFFFE00000, "-2097152.000000"); // -2097152.000000
      convertSigned(32'hCA000000, 64'hFFFFFFFFFFE00000, "-2097152"); // -2097152
      convertSigned(32'hC9FFFFFC, 64'hFFFFFFFFFFE00001, "-2097152.000000"); // -2097152.000000
      convertSigned(32'hC9FFFFF8, 64'hFFFFFFFFFFE00001, "-2097151"); // -2097151
      convertSigned(32'hC9FFFFF4, 64'hFFFFFFFFFFE00002, "-2097150.000000"); // -2097150.000000
      convertSigned(32'hC9800008, 64'hFFFFFFFFFFEFFFFF, "-1048577"); // -1048577
      convertSigned(32'hC9800004, 64'hFFFFFFFFFFF00000, "-1048576.000000"); // -1048576.000000
      convertSigned(32'hC9800000, 64'hFFFFFFFFFFF00000, "-1048576"); // -1048576
      convertSigned(32'hC97FFFF8, 64'hFFFFFFFFFFF00001, "-1048576.000000"); // -1048576.000000
      convertSigned(32'hC97FFFF0, 64'hFFFFFFFFFFF00001, "-1048575"); // -1048575
      convertSigned(32'hC97FFFE8, 64'hFFFFFFFFFFF00002, "-1048574.000000"); // -1048574.000000
      convertSigned(32'hC9000010, 64'hFFFFFFFFFFF7FFFF, "-524289"); // -524289
      convertSigned(32'hC9000008, 64'hFFFFFFFFFFF80000, "-524288.500000"); // -524288.500000
      convertSigned(32'hC9000000, 64'hFFFFFFFFFFF80000, "-524288"); // -524288
      convertSigned(32'hC8FFFFF0, 64'hFFFFFFFFFFF80001, "-524287.500000"); // -524287.500000
      convertSigned(32'hC8FFFFE0, 64'hFFFFFFFFFFF80001, "-524287"); // -524287
      convertSigned(32'hC8FFFFD0, 64'hFFFFFFFFFFF80002, "-524286.500000"); // -524286.500000
      convertSigned(32'hC8800020, 64'hFFFFFFFFFFFBFFFF, "-262145"); // -262145
      convertSigned(32'hC8800010, 64'hFFFFFFFFFFFC0000, "-262144.500000"); // -262144.500000
      convertSigned(32'hC8800000, 64'hFFFFFFFFFFFC0000, "-262144"); // -262144
      convertSigned(32'hC87FFFE0, 64'hFFFFFFFFFFFC0001, "-262143.500000"); // -262143.500000
      convertSigned(32'hC87FFFC0, 64'hFFFFFFFFFFFC0001, "-262143"); // -262143
      convertSigned(32'hC87FFFA0, 64'hFFFFFFFFFFFC0002, "-262142.500000"); // -262142.500000
      convertSigned(32'hC8000040, 64'hFFFFFFFFFFFDFFFF, "-131073"); // -131073
      convertSigned(32'hC8000020, 64'hFFFFFFFFFFFE0000, "-131072.500000"); // -131072.500000
      convertSigned(32'hC8000000, 64'hFFFFFFFFFFFE0000, "-131072"); // -131072
      convertSigned(32'hC7FFFFC0, 64'hFFFFFFFFFFFE0001, "-131071.500000"); // -131071.500000
      convertSigned(32'hC7FFFF80, 64'hFFFFFFFFFFFE0001, "-131071"); // -131071
      convertSigned(32'hC7FFFF40, 64'hFFFFFFFFFFFE0002, "-131070.500000"); // -131070.500000
      convertSigned(32'hC7800080, 64'hFFFFFFFFFFFEFFFF, "-65537"); // -65537
      convertSigned(32'hC7800040, 64'hFFFFFFFFFFFF0000, "-65536.500000"); // -65536.500000
      convertSigned(32'hC7800000, 64'hFFFFFFFFFFFF0000, "-65536"); // -65536
      convertSigned(32'hC77FFF80, 64'hFFFFFFFFFFFF0001, "-65535.500000"); // -65535.500000
      convertSigned(32'hC77FFF00, 64'hFFFFFFFFFFFF0001, "-65535"); // -65535
      convertSigned(32'hC77FFE80, 64'hFFFFFFFFFFFF0002, "-65534.500000"); // -65534.500000
      convertSigned(32'hC7000100, 64'hFFFFFFFFFFFF7FFF, "-32769"); // -32769
      convertSigned(32'hC7000080, 64'hFFFFFFFFFFFF8000, "-32768.500000"); // -32768.500000
      convertSigned(32'hC7000000, 64'hFFFFFFFFFFFF8000, "-32768"); // -32768
      convertSigned(32'hC6FFFF00, 64'hFFFFFFFFFFFF8001, "-32767.500000"); // -32767.500000
      convertSigned(32'hC6FFFE00, 64'hFFFFFFFFFFFF8001, "-32767"); // -32767
      convertSigned(32'hC6FFFD00, 64'hFFFFFFFFFFFF8002, "-32766.500000"); // -32766.500000
      convertSigned(32'hC6800200, 64'hFFFFFFFFFFFFBFFF, "-16385"); // -16385
      convertSigned(32'hC6800100, 64'hFFFFFFFFFFFFC000, "-16384.500000"); // -16384.500000
      convertSigned(32'hC6800000, 64'hFFFFFFFFFFFFC000, "-16384"); // -16384
      convertSigned(32'hC67FFE00, 64'hFFFFFFFFFFFFC001, "-16383.500000"); // -16383.500000
      convertSigned(32'hC67FFC00, 64'hFFFFFFFFFFFFC001, "-16383"); // -16383
      convertSigned(32'hC67FFA00, 64'hFFFFFFFFFFFFC002, "-16382.500000"); // -16382.500000
      convertSigned(32'hC6000400, 64'hFFFFFFFFFFFFDFFF, "-8193"); // -8193
      convertSigned(32'hC6000200, 64'hFFFFFFFFFFFFE000, "-8192.500000"); // -8192.500000
      convertSigned(32'hC6000000, 64'hFFFFFFFFFFFFE000, "-8192"); // -8192
      convertSigned(32'hC5FFFC00, 64'hFFFFFFFFFFFFE001, "-8191.500000"); // -8191.500000
      convertSigned(32'hC5FFF800, 64'hFFFFFFFFFFFFE001, "-8191"); // -8191
      convertSigned(32'hC5FFF400, 64'hFFFFFFFFFFFFE002, "-8190.500000"); // -8190.500000
      convertSigned(32'hC5800800, 64'hFFFFFFFFFFFFEFFF, "-4097"); // -4097
      convertSigned(32'hC5800400, 64'hFFFFFFFFFFFFF000, "-4096.500000"); // -4096.500000
      convertSigned(32'hC5800000, 64'hFFFFFFFFFFFFF000, "-4096"); // -4096
      convertSigned(32'hC57FF800, 64'hFFFFFFFFFFFFF001, "-4095.500000"); // -4095.500000
      convertSigned(32'hC57FF000, 64'hFFFFFFFFFFFFF001, "-4095"); // -4095
      convertSigned(32'hC57FE800, 64'hFFFFFFFFFFFFF002, "-4094.500000"); // -4094.500000
      convertSigned(32'hC5001000, 64'hFFFFFFFFFFFFF7FF, "-2049"); // -2049
      convertSigned(32'hC5000800, 64'hFFFFFFFFFFFFF800, "-2048.500000"); // -2048.500000
      convertSigned(32'hC5000000, 64'hFFFFFFFFFFFFF800, "-2048"); // -2048
      convertSigned(32'hC4FFF000, 64'hFFFFFFFFFFFFF801, "-2047.500000"); // -2047.500000
      convertSigned(32'hC4FFE000, 64'hFFFFFFFFFFFFF801, "-2047"); // -2047
      convertSigned(32'hC4FFD000, 64'hFFFFFFFFFFFFF802, "-2046.500000"); // -2046.500000
      convertSigned(32'hC4802000, 64'hFFFFFFFFFFFFFBFF, "-1025"); // -1025
      convertSigned(32'hC4801000, 64'hFFFFFFFFFFFFFC00, "-1024.500000"); // -1024.500000
      convertSigned(32'hC4800000, 64'hFFFFFFFFFFFFFC00, "-1024"); // -1024
      convertSigned(32'hC47FE000, 64'hFFFFFFFFFFFFFC01, "-1023.500000"); // -1023.500000
      convertSigned(32'hC47FC000, 64'hFFFFFFFFFFFFFC01, "-1023"); // -1023
      convertSigned(32'hC47FA000, 64'hFFFFFFFFFFFFFC02, "-1022.500000"); // -1022.500000
      convertSigned(32'hC4004000, 64'hFFFFFFFFFFFFFDFF, "-513"); // -513
      convertSigned(32'hC4002000, 64'hFFFFFFFFFFFFFE00, "-512.500000"); // -512.500000
      convertSigned(32'hC4000000, 64'hFFFFFFFFFFFFFE00, "-512"); // -512
      convertSigned(32'hC3FFC000, 64'hFFFFFFFFFFFFFE01, "-511.500000"); // -511.500000
      convertSigned(32'hC3FF8000, 64'hFFFFFFFFFFFFFE01, "-511"); // -511
      convertSigned(32'hC3FF4000, 64'hFFFFFFFFFFFFFE02, "-510.500000"); // -510.500000
      convertSigned(32'hC3808000, 64'hFFFFFFFFFFFFFEFF, "-257"); // -257
      convertSigned(32'hC3804000, 64'hFFFFFFFFFFFFFF00, "-256.500000"); // -256.500000
      convertSigned(32'hC3800000, 64'hFFFFFFFFFFFFFF00, "-256"); // -256
      convertSigned(32'hC37F8000, 64'hFFFFFFFFFFFFFF01, "-255.500000"); // -255.500000
      convertSigned(32'hC37F0000, 64'hFFFFFFFFFFFFFF01, "-255"); // -255
      convertSigned(32'hC37E8000, 64'hFFFFFFFFFFFFFF02, "-254.500000"); // -254.500000
      convertSigned(32'hC3010000, 64'hFFFFFFFFFFFFFF7F, "-129"); // -129
      convertSigned(32'hC3008000, 64'hFFFFFFFFFFFFFF80, "-128.500000"); // -128.500000
      convertSigned(32'hC3000000, 64'hFFFFFFFFFFFFFF80, "-128"); // -128
      convertSigned(32'hC2FF0000, 64'hFFFFFFFFFFFFFF81, "-127.500000"); // -127.500000
      convertSigned(32'hC2FE0000, 64'hFFFFFFFFFFFFFF81, "-127"); // -127
      convertSigned(32'hC2FD0000, 64'hFFFFFFFFFFFFFF82, "-126.500000"); // -126.500000
      convertSigned(32'hC2820000, 64'hFFFFFFFFFFFFFFBF, "-65"); // -65
      convertSigned(32'hC2810000, 64'hFFFFFFFFFFFFFFC0, "-64.500000"); // -64.500000
      convertSigned(32'hC2800000, 64'hFFFFFFFFFFFFFFC0, "-64"); // -64
      convertSigned(32'hC27E0000, 64'hFFFFFFFFFFFFFFC1, "-63.500000"); // -63.500000
      convertSigned(32'hC27C0000, 64'hFFFFFFFFFFFFFFC1, "-63"); // -63
      convertSigned(32'hC27A0000, 64'hFFFFFFFFFFFFFFC2, "-62.500000"); // -62.500000
      convertSigned(32'hC2040000, 64'hFFFFFFFFFFFFFFDF, "-33"); // -33
      convertSigned(32'hC2020000, 64'hFFFFFFFFFFFFFFE0, "-32.500000"); // -32.500000
      convertSigned(32'hC2000000, 64'hFFFFFFFFFFFFFFE0, "-32"); // -32
      convertSigned(32'hC1FC0000, 64'hFFFFFFFFFFFFFFE1, "-31.500000"); // -31.500000
      convertSigned(32'hC1F80000, 64'hFFFFFFFFFFFFFFE1, "-31"); // -31
      convertSigned(32'hC1F40000, 64'hFFFFFFFFFFFFFFE2, "-30.500000"); // -30.500000
      convertSigned(32'hC1880000, 64'hFFFFFFFFFFFFFFEF, "-17"); // -17
      convertSigned(32'hC1840000, 64'hFFFFFFFFFFFFFFF0, "-16.500000"); // -16.500000
      convertSigned(32'hC1800000, 64'hFFFFFFFFFFFFFFF0, "-16"); // -16
      convertSigned(32'hC1780000, 64'hFFFFFFFFFFFFFFF1, "-15.500000"); // -15.500000
      convertSigned(32'hC1700000, 64'hFFFFFFFFFFFFFFF1, "-15"); // -15
      convertSigned(32'hC1680000, 64'hFFFFFFFFFFFFFFF2, "-14.500000"); // -14.500000
      convertSigned(32'hC1100000, 64'hFFFFFFFFFFFFFFF7, "-9"); // -9
      convertSigned(32'hC1080000, 64'hFFFFFFFFFFFFFFF8, "-8.500000"); // -8.500000
      convertSigned(32'hC1000000, 64'hFFFFFFFFFFFFFFF8, "-8"); // -8
      convertSigned(32'hC0F00000, 64'hFFFFFFFFFFFFFFF9, "-7.500000"); // -7.500000
      convertSigned(32'hC0E00000, 64'hFFFFFFFFFFFFFFF9, "-7"); // -7
      convertSigned(32'hC0D00000, 64'hFFFFFFFFFFFFFFFA, "-6.500000"); // -6.500000
      convertSigned(32'hC0A00000, 64'hFFFFFFFFFFFFFFFB, "-5"); // -5
      convertSigned(32'hC0900000, 64'hFFFFFFFFFFFFFFFC, "-4.500000"); // -4.500000
      convertSigned(32'hC0800000, 64'hFFFFFFFFFFFFFFFC, "-4"); // -4
      convertSigned(32'hC0600000, 64'hFFFFFFFFFFFFFFFD, "-3.500000"); // -3.500000
      convertSigned(32'hC0400000, 64'hFFFFFFFFFFFFFFFD, "-3"); // -3
      convertSigned(32'hC0200000, 64'hFFFFFFFFFFFFFFFE, "-2.500000"); // -2.500000
      convertSigned(32'hC0000000, 64'hFFFFFFFFFFFFFFFE, "-2"); // -2
      convertSigned(32'hBFC00000, 64'hFFFFFFFFFFFFFFFF, "-1.500000"); // -1.500000
      convertSigned(32'hBF800000, 64'hFFFFFFFFFFFFFFFF, "-1"); // -1
      convertSigned(32'hBF68EFCC, 64'h0000000000000000, "-0.909909"); // -0.909909
      convertSigned(32'hBF143FAC, 64'h0000000000000000, "-0.579097"); // -0.579097
      convertSigned(32'hBF0A2298, 64'h0000000000000000, "-0.539590"); // -0.539590
      convertSigned(32'hBF000000, 64'h0000000000000000, "-0.500000"); // -0.500000
      convertSigned(32'hBECFE64C, 64'h0000000000000000, "-0.406054"); // -0.406054
      convertSigned(32'hBEAA9C2A, 64'h0000000000000000, "-0.333223"); // -0.333223
      convertSigned(32'hBEA44648, 64'h0000000000000000, "-0.320849"); // -0.320849
      convertSigned(32'hBE8A1CBA, 64'h0000000000000000, "-0.269750"); // -0.269750
      convertSigned(32'hBE83870E, 64'h0000000000000000, "-0.256890"); // -0.256890
      convertSigned(32'hBE1906F4, 64'h0000000000000000, "-0.149441"); // -0.149441
      convertSigned(32'h00000000, 64'h0000000000000000, "0"); // 0
      convertSigned(32'h3DF3AB70, 64'h0000000000000000, "0.118979"); // 0.118979
      convertSigned(32'h3E578218, 64'h0000000000000000, "0.210457"); // 0.210457
      convertSigned(32'h3E65B818, 64'h0000000000000000, "0.224335"); // 0.224335
      convertSigned(32'h3E841E7C, 64'h0000000000000000, "0.258045"); // 0.258045
      convertSigned(32'h3E8E39AC, 64'h0000000000000000, "0.277784"); // 0.277784
      convertSigned(32'h3F000000, 64'h0000000000000000, "0.500000"); // 0.500000
      convertSigned(32'h3F25E882, 64'h0000000000000000, "0.648079"); // 0.648079
      convertSigned(32'h3F3441B0, 64'h0000000000000000, "0.704127"); // 0.704127
      convertSigned(32'h3F37E586, 64'h0000000000000000, "0.718346"); // 0.718346
      convertSigned(32'h3F3A5838, 64'h0000000000000000, "0.727909"); // 0.727909
      convertSigned(32'h3F4216A6, 64'h0000000000000000, "0.758158"); // 0.758158
      convertSigned(32'h3F45E488, 64'h0000000000000000, "0.773018"); // 0.773018
      convertSigned(32'h3F800000, 64'h0000000000000001, "1"); // 1
      convertSigned(32'h3FC00000, 64'h0000000000000001, "1.500000"); // 1.500000
      convertSigned(32'h40000000, 64'h0000000000000002, "2"); // 2
      convertSigned(32'h40200000, 64'h0000000000000002, "2.500000"); // 2.500000
      convertSigned(32'h40400000, 64'h0000000000000003, "3"); // 3
      convertSigned(32'h40600000, 64'h0000000000000003, "3.500000"); // 3.500000
      convertSigned(32'h40800000, 64'h0000000000000004, "4"); // 4
      convertSigned(32'h40900000, 64'h0000000000000004, "4.500000"); // 4.500000
      convertSigned(32'h40A00000, 64'h0000000000000005, "5"); // 5
      convertSigned(32'h40B00000, 64'h0000000000000005, "5.500000"); // 5.500000
      convertSigned(32'h40E00000, 64'h0000000000000007, "7"); // 7
      convertSigned(32'h40F00000, 64'h0000000000000007, "7.500000"); // 7.500000
      convertSigned(32'h41000000, 64'h0000000000000008, "8"); // 8
      convertSigned(32'h41080000, 64'h0000000000000008, "8.500000"); // 8.500000
      convertSigned(32'h41100000, 64'h0000000000000009, "9"); // 9
      convertSigned(32'h41180000, 64'h0000000000000009, "9.500000"); // 9.500000
      convertSigned(32'h41700000, 64'h000000000000000F, "15"); // 15
      convertSigned(32'h41780000, 64'h000000000000000F, "15.500000"); // 15.500000
      convertSigned(32'h41800000, 64'h0000000000000010, "16"); // 16
      convertSigned(32'h41840000, 64'h0000000000000010, "16.500000"); // 16.500000
      convertSigned(32'h41880000, 64'h0000000000000011, "17"); // 17
      convertSigned(32'h418C0000, 64'h0000000000000011, "17.500000"); // 17.500000
      convertSigned(32'h41F80000, 64'h000000000000001F, "31"); // 31
      convertSigned(32'h41FC0000, 64'h000000000000001F, "31.500000"); // 31.500000
      convertSigned(32'h42000000, 64'h0000000000000020, "32"); // 32
      convertSigned(32'h42020000, 64'h0000000000000020, "32.500000"); // 32.500000
      convertSigned(32'h42040000, 64'h0000000000000021, "33"); // 33
      convertSigned(32'h42060000, 64'h0000000000000021, "33.500000"); // 33.500000
      convertSigned(32'h427C0000, 64'h000000000000003F, "63"); // 63
      convertSigned(32'h427E0000, 64'h000000000000003F, "63.500000"); // 63.500000
      convertSigned(32'h42800000, 64'h0000000000000040, "64"); // 64
      convertSigned(32'h42810000, 64'h0000000000000040, "64.500000"); // 64.500000
      convertSigned(32'h42820000, 64'h0000000000000041, "65"); // 65
      convertSigned(32'h42830000, 64'h0000000000000041, "65.500000"); // 65.500000
      convertSigned(32'h42FE0000, 64'h000000000000007F, "127"); // 127
      convertSigned(32'h42FF0000, 64'h000000000000007F, "127.500000"); // 127.500000
      convertSigned(32'h43000000, 64'h0000000000000080, "128"); // 128
      convertSigned(32'h43008000, 64'h0000000000000080, "128.500000"); // 128.500000
      convertSigned(32'h43010000, 64'h0000000000000081, "129"); // 129
      convertSigned(32'h43018000, 64'h0000000000000081, "129.500000"); // 129.500000
      convertSigned(32'h437F0000, 64'h00000000000000FF, "255"); // 255
      convertSigned(32'h437F8000, 64'h00000000000000FF, "255.500000"); // 255.500000
      convertSigned(32'h43800000, 64'h0000000000000100, "256"); // 256
      convertSigned(32'h43804000, 64'h0000000000000100, "256.500000"); // 256.500000
      convertSigned(32'h43808000, 64'h0000000000000101, "257"); // 257
      convertSigned(32'h4380C000, 64'h0000000000000101, "257.500000"); // 257.500000
      convertSigned(32'h43FF8000, 64'h00000000000001FF, "511"); // 511
      convertSigned(32'h43FFC000, 64'h00000000000001FF, "511.500000"); // 511.500000
      convertSigned(32'h44000000, 64'h0000000000000200, "512"); // 512
      convertSigned(32'h44002000, 64'h0000000000000200, "512.500000"); // 512.500000
      convertSigned(32'h44004000, 64'h0000000000000201, "513"); // 513
      convertSigned(32'h44006000, 64'h0000000000000201, "513.500000"); // 513.500000
      convertSigned(32'h447FC000, 64'h00000000000003FF, "1023"); // 1023
      convertSigned(32'h447FE000, 64'h00000000000003FF, "1023.500000"); // 1023.500000
      convertSigned(32'h44800000, 64'h0000000000000400, "1024"); // 1024
      convertSigned(32'h44801000, 64'h0000000000000400, "1024.500000"); // 1024.500000
      convertSigned(32'h44802000, 64'h0000000000000401, "1025"); // 1025
      convertSigned(32'h44803000, 64'h0000000000000401, "1025.500000"); // 1025.500000
      convertSigned(32'h44FFE000, 64'h00000000000007FF, "2047"); // 2047
      convertSigned(32'h44FFF000, 64'h00000000000007FF, "2047.500000"); // 2047.500000
      convertSigned(32'h45000000, 64'h0000000000000800, "2048"); // 2048
      convertSigned(32'h45000800, 64'h0000000000000800, "2048.500000"); // 2048.500000
      convertSigned(32'h45001000, 64'h0000000000000801, "2049"); // 2049
      convertSigned(32'h45001800, 64'h0000000000000801, "2049.500000"); // 2049.500000
      convertSigned(32'h457FF000, 64'h0000000000000FFF, "4095"); // 4095
      convertSigned(32'h457FF800, 64'h0000000000000FFF, "4095.500000"); // 4095.500000
      convertSigned(32'h45800000, 64'h0000000000001000, "4096"); // 4096
      convertSigned(32'h45800400, 64'h0000000000001000, "4096.500000"); // 4096.500000
      convertSigned(32'h45800800, 64'h0000000000001001, "4097"); // 4097
      convertSigned(32'h45800C00, 64'h0000000000001001, "4097.500000"); // 4097.500000
      convertSigned(32'h45FFF800, 64'h0000000000001FFF, "8191"); // 8191
      convertSigned(32'h45FFFC00, 64'h0000000000001FFF, "8191.500000"); // 8191.500000
      convertSigned(32'h46000000, 64'h0000000000002000, "8192"); // 8192
      convertSigned(32'h46000200, 64'h0000000000002000, "8192.500000"); // 8192.500000
      convertSigned(32'h46000400, 64'h0000000000002001, "8193"); // 8193
      convertSigned(32'h46000600, 64'h0000000000002001, "8193.500000"); // 8193.500000
      convertSigned(32'h467FFC00, 64'h0000000000003FFF, "16383"); // 16383
      convertSigned(32'h467FFE00, 64'h0000000000003FFF, "16383.500000"); // 16383.500000
      convertSigned(32'h46800000, 64'h0000000000004000, "16384"); // 16384
      convertSigned(32'h46800100, 64'h0000000000004000, "16384.500000"); // 16384.500000
      convertSigned(32'h46800200, 64'h0000000000004001, "16385"); // 16385
      convertSigned(32'h46800300, 64'h0000000000004001, "16385.500000"); // 16385.500000
      convertSigned(32'h46FFFE00, 64'h0000000000007FFF, "32767"); // 32767
      convertSigned(32'h46FFFF00, 64'h0000000000007FFF, "32767.500000"); // 32767.500000
      convertSigned(32'h47000000, 64'h0000000000008000, "32768"); // 32768
      convertSigned(32'h47000080, 64'h0000000000008000, "32768.500000"); // 32768.500000
      convertSigned(32'h47000100, 64'h0000000000008001, "32769"); // 32769
      convertSigned(32'h47000180, 64'h0000000000008001, "32769.500000"); // 32769.500000
      convertSigned(32'h477FFF00, 64'h000000000000FFFF, "65535"); // 65535
      convertSigned(32'h477FFF80, 64'h000000000000FFFF, "65535.500000"); // 65535.500000
      convertSigned(32'h47800000, 64'h0000000000010000, "65536"); // 65536
      convertSigned(32'h47800040, 64'h0000000000010000, "65536.500000"); // 65536.500000
      convertSigned(32'h47800080, 64'h0000000000010001, "65537"); // 65537
      convertSigned(32'h478000C0, 64'h0000000000010001, "65537.500000"); // 65537.500000
      convertSigned(32'h47FFFF80, 64'h000000000001FFFF, "131071"); // 131071
      convertSigned(32'h47FFFFC0, 64'h000000000001FFFF, "131071.500000"); // 131071.500000
      convertSigned(32'h48000000, 64'h0000000000020000, "131072"); // 131072
      convertSigned(32'h48000020, 64'h0000000000020000, "131072.500000"); // 131072.500000
      convertSigned(32'h48000040, 64'h0000000000020001, "131073"); // 131073
      convertSigned(32'h48000060, 64'h0000000000020001, "131073.500000"); // 131073.500000
      convertSigned(32'h487FFFC0, 64'h000000000003FFFF, "262143"); // 262143
      convertSigned(32'h487FFFE0, 64'h000000000003FFFF, "262143.500000"); // 262143.500000
      convertSigned(32'h48800000, 64'h0000000000040000, "262144"); // 262144
      convertSigned(32'h48800010, 64'h0000000000040000, "262144.500000"); // 262144.500000
      convertSigned(32'h48800020, 64'h0000000000040001, "262145"); // 262145
      convertSigned(32'h48800030, 64'h0000000000040001, "262145.500000"); // 262145.500000
      convertSigned(32'h48FFFFE0, 64'h000000000007FFFF, "524287"); // 524287
      convertSigned(32'h48FFFFF0, 64'h000000000007FFFF, "524287.500000"); // 524287.500000
      convertSigned(32'h49000000, 64'h0000000000080000, "524288"); // 524288
      convertSigned(32'h49000008, 64'h0000000000080000, "524288.500000"); // 524288.500000
      convertSigned(32'h49000010, 64'h0000000000080001, "524289"); // 524289
      convertSigned(32'h49000018, 64'h0000000000080001, "524289.500000"); // 524289.500000
      convertSigned(32'h497FFFF0, 64'h00000000000FFFFF, "1048575"); // 1048575
      convertSigned(32'h497FFFF8, 64'h00000000000FFFFF, "1048576.000000"); // 1048576.000000
      convertSigned(32'h49800000, 64'h0000000000100000, "1048576"); // 1048576
      convertSigned(32'h49800004, 64'h0000000000100000, "1048576.000000"); // 1048576.000000
      convertSigned(32'h49800008, 64'h0000000000100001, "1048577"); // 1048577
      convertSigned(32'h4980000C, 64'h0000000000100001, "1048578.000000"); // 1048578.000000
      convertSigned(32'h49FFFFF8, 64'h00000000001FFFFF, "2097151"); // 2097151
      convertSigned(32'h49FFFFFC, 64'h00000000001FFFFF, "2097152.000000"); // 2097152.000000
      convertSigned(32'h4A000000, 64'h0000000000200000, "2097152"); // 2097152
      convertSigned(32'h4A000002, 64'h0000000000200000, "2097152.000000"); // 2097152.000000
      convertSigned(32'h4A000004, 64'h0000000000200001, "2097153"); // 2097153
      convertSigned(32'h4A000006, 64'h0000000000200001, "2097154.000000"); // 2097154.000000
      convertSigned(32'h4A7FFFFC, 64'h00000000003FFFFF, "4194303"); // 4194303
      convertSigned(32'h4A7FFFFE, 64'h00000000003FFFFF, "4194304.000000"); // 4194304.000000
      convertSigned(32'h4A800000, 64'h0000000000400000, "4194304"); // 4194304
      convertSigned(32'h4A800001, 64'h0000000000400000, "4194304.000000"); // 4194304.000000
      convertSigned(32'h4A800002, 64'h0000000000400001, "4194305"); // 4194305
      convertSigned(32'h4A800003, 64'h0000000000400001, "4194306.000000"); // 4194306.000000
      convertSigned(32'h4AFFFFFE, 64'h00000000007FFFFF, "8388607"); // 8388607
      convertSigned(32'h4AFFFFFF, 64'h00000000007FFFFF, "8388608.000000"); // 8388608.000000
      convertSigned(32'h4B000000, 64'h0000000000800000, "8388608.000000"); // 8388608.000000
      convertSigned(32'h4B000001, 64'h0000000000800001, "8388609"); // 8388609
      convertSigned(32'h4B000002, 64'h0000000000800002, "8388610.000000"); // 8388610.000000
      convertSigned(32'h4B800000, 64'h0000000001000000, "16777220.000000"); // 16777220.000000
      convertSigned(32'h4B800001, 64'h0000000001000002, "16777220.000000"); // 16777220.000000
      convertSigned(32'h4B800002, 64'h0000000001000004, "16777220.000000"); // 16777220.000000
      convertSigned(32'h4C000000, 64'h0000000002000000, "33554430.000000"); // 33554430.000000
      convertSigned(32'h4C000001, 64'h0000000002000004, "33554440.000000"); // 33554440.000000
      convertSigned(32'h4C000002, 64'h0000000002000008, "33554440.000000"); // 33554440.000000
      convertSigned(32'h4C800000, 64'h0000000004000000, "67108860.000000"); // 67108860.000000
      convertSigned(32'h4C800001, 64'h0000000004000008, "67108870.000000"); // 67108870.000000
      convertSigned(32'h4C800002, 64'h0000000004000010, "67108880.000000"); // 67108880.000000
      convertSigned(32'h4D000000, 64'h0000000008000000, "134217700.000000"); // 134217700.000000
      convertSigned(32'h4D000001, 64'h0000000008000010, "134217700.000000"); // 134217700.000000
      convertSigned(32'h4D000002, 64'h0000000008000020, "134217800.000000"); // 134217800.000000
      convertSigned(32'h4D800000, 64'h0000000010000000, "268435500.000000"); // 268435500.000000
      convertSigned(32'h4D800001, 64'h0000000010000020, "268435500.000000"); // 268435500.000000
      convertSigned(32'h4D800002, 64'h0000000010000040, "268435500.000000"); // 268435500.000000
      convertSigned(32'h4E000000, 64'h0000000020000000, "536870900.000000"); // 536870900.000000
      convertSigned(32'h4E000001, 64'h0000000020000040, "536871000.000000"); // 536871000.000000
      convertSigned(32'h4E000002, 64'h0000000020000080, "536871000.000000"); // 536871000.000000
      convertSigned(32'h4E800000, 64'h0000000040000000, "1073742000.000000"); // 1073742000.000000
      convertSigned(32'h4E800001, 64'h0000000040000080, "1073742000.000000"); // 1073742000.000000
      convertSigned(32'h4E800002, 64'h0000000040000100, "1073742000.000000"); // 1073742000.000000
      convertSigned(32'h4F000000, 64'h0000000080000000, "2147484000.000000"); // 2147484000.000000
      convertSigned(32'h4F000001, 64'h0000000080000100, "2147484000.000000"); // 2147484000.000000
      convertSigned(32'h4F000002, 64'h0000000080000200, "2147484000.000000"); // 2147484000.000000
      convertSigned(32'h4F800000, 64'h0000000100000000, "4294967000.000000"); // 4294967000.000000
      convertSigned(32'h4F800001, 64'h0000000100000200, "4294968000.000000"); // 4294968000.000000
      convertSigned(32'h4F800002, 64'h0000000100000400, "4294968000.000000"); // 4294968000.000000
      convertSigned(32'h50000000, 64'h0000000200000000, "8589935000.000000"); // 8589935000.000000
      convertSigned(32'h50000001, 64'h0000000200000400, "8589936000.000000"); // 8589936000.000000
      convertSigned(32'h50000002, 64'h0000000200000800, "8589937000.000000"); // 8589937000.000000
      convertSigned(32'h50800000, 64'h0000000400000000, "17179870000.000000"); // 17179870000.000000
      convertSigned(32'h50800001, 64'h0000000400000800, "17179870000.000000"); // 17179870000.000000
      convertSigned(32'h50800002, 64'h0000000400001000, "17179870000.000000"); // 17179870000.000000
      convertSigned(32'h51000000, 64'h0000000800000000, "34359740000.000000"); // 34359740000.000000
      convertSigned(32'h51000001, 64'h0000000800001000, "34359740000.000000"); // 34359740000.000000
      convertSigned(32'h51000002, 64'h0000000800002000, "34359750000.000000"); // 34359750000.000000
      convertSigned(32'h51800000, 64'h0000001000000000, "68719480000.000000"); // 68719480000.000000
      convertSigned(32'h51800001, 64'h0000001000002000, "68719480000.000000"); // 68719480000.000000
      convertSigned(32'h51800002, 64'h0000001000004000, "68719490000.000000"); // 68719490000.000000
      convertSigned(32'h52000000, 64'h0000002000000000, "137439000000.000000"); // 137439000000.000000
      convertSigned(32'h52000001, 64'h0000002000004000, "137439000000.000000"); // 137439000000.000000
      convertSigned(32'h52000002, 64'h0000002000008000, "137439000000.000000"); // 137439000000.000000
      convertSigned(32'h52800000, 64'h0000004000000000, "274877900000.000000"); // 274877900000.000000
      convertSigned(32'h52800001, 64'h0000004000008000, "274877900000.000000"); // 274877900000.000000
      convertSigned(32'h52800002, 64'h0000004000010000, "274878000000.000000"); // 274878000000.000000
      convertSigned(32'h53000000, 64'h0000008000000000, "549755800000.000000"); // 549755800000.000000
      convertSigned(32'h53000001, 64'h0000008000010000, "549755900000.000000"); // 549755900000.000000
      convertSigned(32'h53000002, 64'h0000008000020000, "549755900000.000000"); // 549755900000.000000
      convertSigned(32'h53800000, 64'h0000010000000000, "1099512000000.000000"); // 1099512000000.000000
      convertSigned(32'h53800001, 64'h0000010000020000, "1099512000000.000000"); // 1099512000000.000000
      convertSigned(32'h53800002, 64'h0000010000040000, "1099512000000.000000"); // 1099512000000.000000
      convertSigned(32'h54000000, 64'h0000020000000000, "2199023000000.000000"); // 2199023000000.000000
      convertSigned(32'h54000001, 64'h0000020000040000, "2199024000000.000000"); // 2199024000000.000000
      convertSigned(32'h54000002, 64'h0000020000080000, "2199024000000.000000"); // 2199024000000.000000
      convertSigned(32'h54800000, 64'h0000040000000000, "4398047000000.000000"); // 4398047000000.000000
      convertSigned(32'h54800001, 64'h0000040000080000, "4398047000000.000000"); // 4398047000000.000000
      convertSigned(32'h54800002, 64'h0000040000100000, "4398048000000.000000"); // 4398048000000.000000
      convertSigned(32'h55000000, 64'h0000080000000000, "8796093000000.000000"); // 8796093000000.000000
      convertSigned(32'h55000001, 64'h0000080000100000, "8796094000000.000000"); // 8796094000000.000000
      convertSigned(32'h55000002, 64'h0000080000200000, "8796095000000.000000"); // 8796095000000.000000
      convertSigned(32'h55800000, 64'h0000100000000000, "17592190000000.000000"); // 17592190000000.000000
      convertSigned(32'h55800001, 64'h0000100000200000, "17592190000000.000000"); // 17592190000000.000000
      convertSigned(32'h55800002, 64'h0000100000400000, "17592190000000.000000"); // 17592190000000.000000
      convertSigned(32'h56000000, 64'h0000200000000000, "35184370000000.000000"); // 35184370000000.000000
      convertSigned(32'h56000001, 64'h0000200000400000, "35184380000000.000000"); // 35184380000000.000000
      convertSigned(32'h56000002, 64'h0000200000800000, "35184380000000.000000"); // 35184380000000.000000
      convertSigned(32'h56800000, 64'h0000400000000000, "70368740000000.000000"); // 70368740000000.000000
      convertSigned(32'h56800001, 64'h0000400000800000, "70368750000000.000000"); // 70368750000000.000000
      convertSigned(32'h56800002, 64'h0000400001000000, "70368760000000.000000"); // 70368760000000.000000
      convertSigned(32'h57000000, 64'h0000800000000000, "140737500000000.000000"); // 140737500000000.000000
      convertSigned(32'h57000001, 64'h0000800001000000, "140737500000000.000000"); // 140737500000000.000000
      convertSigned(32'h57000002, 64'h0000800002000000, "140737500000000.000000"); // 140737500000000.000000
      convertSigned(32'h57800000, 64'h0001000000000000, "281475000000000.000000"); // 281475000000000.000000
      convertSigned(32'h57800001, 64'h0001000002000000, "281475000000000.000000"); // 281475000000000.000000
      convertSigned(32'h57800002, 64'h0001000004000000, "281475000000000.000000"); // 281475000000000.000000
      convertSigned(32'h58000000, 64'h0002000000000000, "562950000000000.000000"); // 562950000000000.000000
      convertSigned(32'h58000001, 64'h0002000004000000, "562950000000000.000000"); // 562950000000000.000000
      convertSigned(32'h58000002, 64'h0002000008000000, "562950100000000.000000"); // 562950100000000.000000
      convertSigned(32'h58800000, 64'h0004000000000000, "1125900000000000.000000"); // 1125900000000000.000000
      convertSigned(32'h58800001, 64'h0004000008000000, "1125900000000000.000000"); // 1125900000000000.000000
      convertSigned(32'h58800002, 64'h0004000010000000, "1125900000000000.000000"); // 1125900000000000.000000
      convertSigned(32'h59000000, 64'h0008000000000000, "2251800000000000.000000"); // 2251800000000000.000000
      convertSigned(32'h59000001, 64'h0008000010000000, "2251800000000000.000000"); // 2251800000000000.000000
      convertSigned(32'h59000002, 64'h0008000020000000, "2251800000000000.000000"); // 2251800000000000.000000
      convertSigned(32'h59800000, 64'h0010000000000000, "4503600000000000.000000"); // 4503600000000000.000000
      convertSigned(32'h59800001, 64'h0010000020000000, "4503600000000000.000000"); // 4503600000000000.000000
      convertSigned(32'h59800002, 64'h0010000040000000, "4503601000000000.000000"); // 4503601000000000.000000
      convertSigned(32'h5A000000, 64'h0020000000000000, "9007199000000000.000000"); // 9007199000000000.000000
      convertSigned(32'h5A000001, 64'h0020000040000000, "9007200000000000.000000"); // 9007200000000000.000000
      convertSigned(32'h5A000002, 64'h0020000080000000, "9007201000000000.000000"); // 9007201000000000.000000
      convertSigned(32'h5A800000, 64'h0040000000000000, "18014400000000000.000000"); // 18014400000000000.000000
      convertSigned(32'h5A800001, 64'h0040000080000000, "18014400000000000.000000"); // 18014400000000000.000000
      convertSigned(32'h5A800002, 64'h0040000100000000, "18014400000000000.000000"); // 18014400000000000.000000
      convertSigned(32'h5B000000, 64'h0080000000000000, "36028800000000000.000000"); // 36028800000000000.000000
      convertSigned(32'h5B000001, 64'h0080000100000000, "36028800000000000.000000"); // 36028800000000000.000000
      convertSigned(32'h5B000002, 64'h0080000200000000, "36028810000000000.000000"); // 36028810000000000.000000
      convertSigned(32'h5B800000, 64'h0100000000000000, "72057590000000000.000000"); // 72057590000000000.000000
      convertSigned(32'h5B800001, 64'h0100000200000000, "72057600000000000.000000"); // 72057600000000000.000000
      convertSigned(32'h5B800002, 64'h0100000400000000, "72057610000000000.000000"); // 72057610000000000.000000
      convertSigned(32'h5C000000, 64'h0200000000000000, "144115200000000000.000000"); // 144115200000000000.000000
      convertSigned(32'h5C000001, 64'h0200000400000000, "144115200000000000.000000"); // 144115200000000000.000000
      convertSigned(32'h5C000002, 64'h0200000800000000, "144115200000000000.000000"); // 144115200000000000.000000
      convertSigned(32'h5C800000, 64'h0400000000000000, "288230400000000000.000000"); // 288230400000000000.000000
      convertSigned(32'h5C800001, 64'h0400000800000000, "288230400000000000.000000"); // 288230400000000000.000000
      convertSigned(32'h5C800002, 64'h0400001000000000, "288230400000000000.000000"); // 288230400000000000.000000
      convertSigned(32'h5D000000, 64'h0800000000000000, "576460800000000000.000000"); // 576460800000000000.000000
      convertSigned(32'h5D000001, 64'h0800001000000000, "576460800000000000.000000"); // 576460800000000000.000000
      convertSigned(32'h5D000002, 64'h0800002000000000, "576460900000000000.000000"); // 576460900000000000.000000
      convertSigned(32'h5D800000, 64'h1000000000000000, "1152922000000000000.000000"); // 1152922000000000000.000000
      convertSigned(32'h5D800001, 64'h1000002000000000, "1152922000000000000.000000"); // 1152922000000000000.000000
      convertSigned(32'h5D800002, 64'h1000004000000000, "1152922000000000000.000000"); // 1152922000000000000.000000
      convertSigned(32'h5E000000, 64'h2000000000000000, "2305843000000000000.000000"); // 2305843000000000000.000000
      convertSigned(32'h5E000001, 64'h2000004000000000, "2305843000000000000.000000"); // 2305843000000000000.000000
      convertSigned(32'h5E000002, 64'h2000008000000000, "2305844000000000000.000000"); // 2305844000000000000.000000
      convertSigned(32'h5E800000, 64'h4000000000000000, "4611686000000000000.000000"); // 4611686000000000000.000000
      convertSigned(32'h5E800001, 64'h4000008000000000, "4611687000000000000.000000"); // 4611687000000000000.000000
      convertSigned(32'h5E800002, 64'h4000010000000000, "4611687000000000000.000000"); // 4611687000000000000.000000
      convertSigned(32'h7F800000, 64'h8000000000000000, "Pos Inf"); // Pos Inf
      
    end
    `uvm_info("LABEL", "Finished run phase.", UVM_HIGH);
    phase.drop_objection(this);
  endtask: run_phase
  
endclass

//-----------
// module top
//-----------
module top;

  bit clk;
  env environment;
  FloatToInt dut(.clk (clk));

  initial begin
    environment = new("env");
    // Put the interface into the resource database.
    uvm_resource_db#(virtual FloatToInt_IF)::set("env",
      "FloatToInt_IF", dut.FloatToInt_IF0);
    clk = 0;
    run_test();
  end
  
  initial begin
    forever begin
      #(50) clk = ~clk;
    end
  end
  
  initial begin
    // Dump waves
    $dumpvars(0, top);
  end
  
endmodule