/*
 *  64 bit integer to float converter
 *
 *  Copyright (C) 2019  Evgeny Muryshkin <evmuryshkin@gmail.com>
 *
 *  Part of Quokka FPGA toolkit
 *  https://github.com/EvgenyMuryshkin/QuokkaEvaluation
 *
 *  Permission to use, copy, modify, and/or distribute this software for any
 *  purpose with or without fee is hereby granted, provided that the above
 *  copyright notice and this permission notice appear in all copies.
 *
 *  THE SOFTWARE IS PROVIDED "AS IS" AND THE AUTHOR DISCLAIMS ALL WARRANTIES
 *  WITH REGARD TO THIS SOFTWARE INCLUDING ALL IMPLIED WARRANTIES OF
 *  MERCHANTABILITY AND FITNESS. IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR
 *  ANY SPECIAL, DIRECT, INDIRECT, OR CONSEQUENTIAL DAMAGES OR ANY DAMAGES
 *  WHATSOEVER RESULTING FROM LOSS OF USE, DATA OR PROFITS, WHETHER IN AN
 *  ACTION OF CONTRACT, NEGLIGENCE OR OTHER TORTIOUS ACTION, ARISING OUT OF
 *  OR IN CONNECTION WITH THE USE OR PERFORMANCE OF THIS SOFTWARE.
 */
import uvm_pkg::*;
`include "uvm_macros.svh"

//---------------------------------------
// Interface for the IntToFloat DUT
//---------------------------------------
interface IntToFloat_IF(
	input bit clk,
  	input inTrigger,
  	input inIsSigned,
	input [63:0] inData,
	input [31:0] outData,
	input outReady
);

  clocking cb @(posedge clk);
    output     inTrigger;
    output     inIsSigned;
    output     inData;
    input    outData;
    input    outReady;
  endclocking // cb

endinterface: IntToFloat_IF

//---------------
// Interface bind
//---------------
bind IntToFloat IntToFloat_IF IntToFloat_IF0(
  .clk(clk),
  .inTrigger(inTrigger),
  .inIsSigned(inIsSigned),
  .inData(inData),
  .outData(outData),
  .outReady(outReady)
);

//----------------
// environment env
//----------------
class env extends uvm_env;

  virtual IntToFloat_IF m_if;

  function new(string name, uvm_component parent = null);
    super.new(name, parent);
  endfunction
  
  function void connect_phase(uvm_phase phase);
    `uvm_info("LABEL", "Started connect phase.", UVM_HIGH);
    // Get the interface from the resource database.
    assert(uvm_resource_db#(virtual IntToFloat_IF)::read_by_name(
      get_full_name(), "IntToFloat_IF", m_if));
    `uvm_info("LABEL", "Finished connect phase.", UVM_HIGH);
  endfunction: connect_phase

  task fullCycle();
    begin
      repeat(2) @(m_if.cb);
    end
  endtask
  
  task convertSigned(longint value, int unsigned expected);
    begin
      m_if.cb.inData <= value;
      m_if.cb.inIsSigned <= 1;
      m_if.cb.inTrigger <= 1;
      fullCycle();
      
      m_if.cb.inTrigger <= 0;
      repeat(64) fullCycle();

      `uvm_info("RESULT", $sformatf("%0d[%0x] = %0x", value, expected, m_if.cb.outData), UVM_LOW);
      if (m_if.cb.outReady != 1)
        `uvm_error("outReady", "Did not finish convertion");
      
      if (m_if.cb.outData != expected)
        `uvm_error("outData", "Result did not match");

    end
  endtask
  
  task run_phase(uvm_phase phase);
    phase.raise_objection(this);
    `uvm_info("LABEL", "Started run phase.", UVM_HIGH);
    begin
      @(m_if.cb);
     
      // incremental bits signed test cases
      convertSigned(64'h0000000000000000, 32'h00000000); // 0
      convertSigned(64'h0000000000000000, 32'h00000000); // 0
      convertSigned(64'h0000000000000001, 32'h3F800000); // 1
      convertSigned(64'hFFFFFFFFFFFFFFFF, 32'hBF800000); // -1
      convertSigned(64'h0000000000000002, 32'h40000000); // 2
      convertSigned(64'hFFFFFFFFFFFFFFFE, 32'hC0000000); // -2
      convertSigned(64'h0000000000000001, 32'h3F800000); // 1
      convertSigned(64'hFFFFFFFFFFFFFFFF, 32'hBF800000); // -1
      convertSigned(64'h0000000000000002, 32'h40000000); // 2
      convertSigned(64'hFFFFFFFFFFFFFFFE, 32'hC0000000); // -2
      convertSigned(64'h0000000000000003, 32'h40400000); // 3
      convertSigned(64'hFFFFFFFFFFFFFFFD, 32'hC0400000); // -3
      convertSigned(64'h0000000000000003, 32'h40400000); // 3
      convertSigned(64'hFFFFFFFFFFFFFFFD, 32'hC0400000); // -3
      convertSigned(64'h0000000000000004, 32'h40800000); // 4
      convertSigned(64'hFFFFFFFFFFFFFFFC, 32'hC0800000); // -4
      convertSigned(64'h0000000000000005, 32'h40A00000); // 5
      convertSigned(64'hFFFFFFFFFFFFFFFB, 32'hC0A00000); // -5
      convertSigned(64'h0000000000000007, 32'h40E00000); // 7
      convertSigned(64'hFFFFFFFFFFFFFFF9, 32'hC0E00000); // -7
      convertSigned(64'h0000000000000008, 32'h41000000); // 8
      convertSigned(64'hFFFFFFFFFFFFFFF8, 32'hC1000000); // -8
      convertSigned(64'h0000000000000009, 32'h41100000); // 9
      convertSigned(64'hFFFFFFFFFFFFFFF7, 32'hC1100000); // -9
      convertSigned(64'h000000000000000F, 32'h41700000); // 15
      convertSigned(64'hFFFFFFFFFFFFFFF1, 32'hC1700000); // -15
      convertSigned(64'h0000000000000010, 32'h41800000); // 16
      convertSigned(64'hFFFFFFFFFFFFFFF0, 32'hC1800000); // -16
      convertSigned(64'h0000000000000011, 32'h41880000); // 17
      convertSigned(64'hFFFFFFFFFFFFFFEF, 32'hC1880000); // -17
      convertSigned(64'h000000000000001F, 32'h41F80000); // 31
      convertSigned(64'hFFFFFFFFFFFFFFE1, 32'hC1F80000); // -31
      convertSigned(64'h0000000000000020, 32'h42000000); // 32
      convertSigned(64'hFFFFFFFFFFFFFFE0, 32'hC2000000); // -32
      convertSigned(64'h0000000000000021, 32'h42040000); // 33
      convertSigned(64'hFFFFFFFFFFFFFFDF, 32'hC2040000); // -33
      convertSigned(64'h000000000000003F, 32'h427C0000); // 63
      convertSigned(64'hFFFFFFFFFFFFFFC1, 32'hC27C0000); // -63
      convertSigned(64'h0000000000000040, 32'h42800000); // 64
      convertSigned(64'hFFFFFFFFFFFFFFC0, 32'hC2800000); // -64
      convertSigned(64'h0000000000000041, 32'h42820000); // 65
      convertSigned(64'hFFFFFFFFFFFFFFBF, 32'hC2820000); // -65
      convertSigned(64'h000000000000007F, 32'h42FE0000); // 127
      convertSigned(64'hFFFFFFFFFFFFFF81, 32'hC2FE0000); // -127
      convertSigned(64'h0000000000000080, 32'h43000000); // 128
      convertSigned(64'hFFFFFFFFFFFFFF80, 32'hC3000000); // -128
      convertSigned(64'h0000000000000081, 32'h43010000); // 129
      convertSigned(64'hFFFFFFFFFFFFFF7F, 32'hC3010000); // -129
      convertSigned(64'h00000000000000FF, 32'h437F0000); // 255
      convertSigned(64'hFFFFFFFFFFFFFF01, 32'hC37F0000); // -255
      convertSigned(64'h0000000000000100, 32'h43800000); // 256
      convertSigned(64'hFFFFFFFFFFFFFF00, 32'hC3800000); // -256
      convertSigned(64'h0000000000000101, 32'h43808000); // 257
      convertSigned(64'hFFFFFFFFFFFFFEFF, 32'hC3808000); // -257
      convertSigned(64'h00000000000001FF, 32'h43FF8000); // 511
      convertSigned(64'hFFFFFFFFFFFFFE01, 32'hC3FF8000); // -511
      convertSigned(64'h0000000000000200, 32'h44000000); // 512
      convertSigned(64'hFFFFFFFFFFFFFE00, 32'hC4000000); // -512
      convertSigned(64'h0000000000000201, 32'h44004000); // 513
      convertSigned(64'hFFFFFFFFFFFFFDFF, 32'hC4004000); // -513
      convertSigned(64'h00000000000003FF, 32'h447FC000); // 1023
      convertSigned(64'hFFFFFFFFFFFFFC01, 32'hC47FC000); // -1023
      convertSigned(64'h0000000000000400, 32'h44800000); // 1024
      convertSigned(64'hFFFFFFFFFFFFFC00, 32'hC4800000); // -1024
      convertSigned(64'h0000000000000401, 32'h44802000); // 1025
      convertSigned(64'hFFFFFFFFFFFFFBFF, 32'hC4802000); // -1025
      convertSigned(64'h00000000000007FF, 32'h44FFE000); // 2047
      convertSigned(64'hFFFFFFFFFFFFF801, 32'hC4FFE000); // -2047
      convertSigned(64'h0000000000000800, 32'h45000000); // 2048
      convertSigned(64'hFFFFFFFFFFFFF800, 32'hC5000000); // -2048
      convertSigned(64'h0000000000000801, 32'h45001000); // 2049
      convertSigned(64'hFFFFFFFFFFFFF7FF, 32'hC5001000); // -2049
      convertSigned(64'h0000000000000FFF, 32'h457FF000); // 4095
      convertSigned(64'hFFFFFFFFFFFFF001, 32'hC57FF000); // -4095
      convertSigned(64'h0000000000001000, 32'h45800000); // 4096
      convertSigned(64'hFFFFFFFFFFFFF000, 32'hC5800000); // -4096
      convertSigned(64'h0000000000001001, 32'h45800800); // 4097
      convertSigned(64'hFFFFFFFFFFFFEFFF, 32'hC5800800); // -4097
      convertSigned(64'h0000000000001FFF, 32'h45FFF800); // 8191
      convertSigned(64'hFFFFFFFFFFFFE001, 32'hC5FFF800); // -8191
      convertSigned(64'h0000000000002000, 32'h46000000); // 8192
      convertSigned(64'hFFFFFFFFFFFFE000, 32'hC6000000); // -8192
      convertSigned(64'h0000000000002001, 32'h46000400); // 8193
      convertSigned(64'hFFFFFFFFFFFFDFFF, 32'hC6000400); // -8193
      convertSigned(64'h0000000000003FFF, 32'h467FFC00); // 16383
      convertSigned(64'hFFFFFFFFFFFFC001, 32'hC67FFC00); // -16383
      convertSigned(64'h0000000000004000, 32'h46800000); // 16384
      convertSigned(64'hFFFFFFFFFFFFC000, 32'hC6800000); // -16384
      convertSigned(64'h0000000000004001, 32'h46800200); // 16385
      convertSigned(64'hFFFFFFFFFFFFBFFF, 32'hC6800200); // -16385
      convertSigned(64'h0000000000007FFF, 32'h46FFFE00); // 32767
      convertSigned(64'hFFFFFFFFFFFF8001, 32'hC6FFFE00); // -32767
      convertSigned(64'h0000000000008000, 32'h47000000); // 32768
      convertSigned(64'hFFFFFFFFFFFF8000, 32'hC7000000); // -32768
      convertSigned(64'h0000000000008001, 32'h47000100); // 32769
      convertSigned(64'hFFFFFFFFFFFF7FFF, 32'hC7000100); // -32769
      convertSigned(64'h000000000000FFFF, 32'h477FFF00); // 65535
      convertSigned(64'hFFFFFFFFFFFF0001, 32'hC77FFF00); // -65535
      convertSigned(64'h0000000000010000, 32'h47800000); // 65536
      convertSigned(64'hFFFFFFFFFFFF0000, 32'hC7800000); // -65536
      convertSigned(64'h0000000000010001, 32'h47800080); // 65537
      convertSigned(64'hFFFFFFFFFFFEFFFF, 32'hC7800080); // -65537
      convertSigned(64'h000000000001FFFF, 32'h47FFFF80); // 131071
      convertSigned(64'hFFFFFFFFFFFE0001, 32'hC7FFFF80); // -131071
      convertSigned(64'h0000000000020000, 32'h48000000); // 131072
      convertSigned(64'hFFFFFFFFFFFE0000, 32'hC8000000); // -131072
      convertSigned(64'h0000000000020001, 32'h48000040); // 131073
      convertSigned(64'hFFFFFFFFFFFDFFFF, 32'hC8000040); // -131073
      convertSigned(64'h000000000003FFFF, 32'h487FFFC0); // 262143
      convertSigned(64'hFFFFFFFFFFFC0001, 32'hC87FFFC0); // -262143
      convertSigned(64'h0000000000040000, 32'h48800000); // 262144
      convertSigned(64'hFFFFFFFFFFFC0000, 32'hC8800000); // -262144
      convertSigned(64'h0000000000040001, 32'h48800020); // 262145
      convertSigned(64'hFFFFFFFFFFFBFFFF, 32'hC8800020); // -262145
      convertSigned(64'h000000000007FFFF, 32'h48FFFFE0); // 524287
      convertSigned(64'hFFFFFFFFFFF80001, 32'hC8FFFFE0); // -524287
      convertSigned(64'h0000000000080000, 32'h49000000); // 524288
      convertSigned(64'hFFFFFFFFFFF80000, 32'hC9000000); // -524288
      convertSigned(64'h0000000000080001, 32'h49000010); // 524289
      convertSigned(64'hFFFFFFFFFFF7FFFF, 32'hC9000010); // -524289
      convertSigned(64'h00000000000FFFFF, 32'h497FFFF0); // 1048575
      convertSigned(64'hFFFFFFFFFFF00001, 32'hC97FFFF0); // -1048575
      convertSigned(64'h0000000000100000, 32'h49800000); // 1048576
      convertSigned(64'hFFFFFFFFFFF00000, 32'hC9800000); // -1048576
      convertSigned(64'h0000000000100001, 32'h49800008); // 1048577
      convertSigned(64'hFFFFFFFFFFEFFFFF, 32'hC9800008); // -1048577
      convertSigned(64'h00000000001FFFFF, 32'h49FFFFF8); // 2097151
      convertSigned(64'hFFFFFFFFFFE00001, 32'hC9FFFFF8); // -2097151
      convertSigned(64'h0000000000200000, 32'h4A000000); // 2097152
      convertSigned(64'hFFFFFFFFFFE00000, 32'hCA000000); // -2097152
      convertSigned(64'h0000000000200001, 32'h4A000004); // 2097153
      convertSigned(64'hFFFFFFFFFFDFFFFF, 32'hCA000004); // -2097153
      convertSigned(64'h00000000003FFFFF, 32'h4A7FFFFC); // 4194303
      convertSigned(64'hFFFFFFFFFFC00001, 32'hCA7FFFFC); // -4194303
      convertSigned(64'h0000000000400000, 32'h4A800000); // 4194304
      convertSigned(64'hFFFFFFFFFFC00000, 32'hCA800000); // -4194304
      convertSigned(64'h0000000000400001, 32'h4A800002); // 4194305
      convertSigned(64'hFFFFFFFFFFBFFFFF, 32'hCA800002); // -4194305
      convertSigned(64'h00000000007FFFFF, 32'h4AFFFFFE); // 8388607
      convertSigned(64'hFFFFFFFFFF800001, 32'hCAFFFFFE); // -8388607
      convertSigned(64'h0000000000800000, 32'h4B000000); // 8388608
      convertSigned(64'hFFFFFFFFFF800000, 32'hCB000000); // -8388608
      convertSigned(64'h0000000000800001, 32'h4B000001); // 8388609
      convertSigned(64'hFFFFFFFFFF7FFFFF, 32'hCB000001); // -8388609
      convertSigned(64'h0000000001000000, 32'h4B800000); // 16777216
      convertSigned(64'hFFFFFFFFFF000000, 32'hCB800000); // -16777216
      convertSigned(64'h0000000001000001, 32'h4B800000); // 16777217
      convertSigned(64'hFFFFFFFFFEFFFFFF, 32'hCB800000); // -16777217
      convertSigned(64'h0000000001000002, 32'h4B800001); // 16777218
      convertSigned(64'hFFFFFFFFFEFFFFFE, 32'hCB800001); // -16777218
      convertSigned(64'h0000000001000002, 32'h4B800001); // 16777218
      convertSigned(64'hFFFFFFFFFEFFFFFE, 32'hCB800001); // -16777218
      convertSigned(64'h0000000001000003, 32'h4B800002); // 16777219
      convertSigned(64'hFFFFFFFFFEFFFFFD, 32'hCB800002); // -16777219
      convertSigned(64'h0000000001000004, 32'h4B800002); // 16777220
      convertSigned(64'hFFFFFFFFFEFFFFFC, 32'hCB800002); // -16777220
      convertSigned(64'h0000000002000001, 32'h4C000000); // 33554433
      convertSigned(64'hFFFFFFFFFDFFFFFF, 32'hCC000000); // -33554433
      convertSigned(64'h0000000002000002, 32'h4C000000); // 33554434
      convertSigned(64'hFFFFFFFFFDFFFFFE, 32'hCC000000); // -33554434
      convertSigned(64'h0000000002000003, 32'h4C000001); // 33554435
      convertSigned(64'hFFFFFFFFFDFFFFFD, 32'hCC000001); // -33554435
      convertSigned(64'h0000000002000005, 32'h4C000001); // 33554437
      convertSigned(64'hFFFFFFFFFDFFFFFB, 32'hCC000001); // -33554437
      convertSigned(64'h0000000002000006, 32'h4C000002); // 33554438
      convertSigned(64'hFFFFFFFFFDFFFFFA, 32'hCC000002); // -33554438
      convertSigned(64'h0000000002000007, 32'h4C000002); // 33554439
      convertSigned(64'hFFFFFFFFFDFFFFF9, 32'hCC000002); // -33554439
      convertSigned(64'h0000000004000003, 32'h4C800000); // 67108867
      convertSigned(64'hFFFFFFFFFBFFFFFD, 32'hCC800000); // -67108867
      convertSigned(64'h0000000004000004, 32'h4C800000); // 67108868
      convertSigned(64'hFFFFFFFFFBFFFFFC, 32'hCC800000); // -67108868
      convertSigned(64'h0000000004000005, 32'h4C800001); // 67108869
      convertSigned(64'hFFFFFFFFFBFFFFFB, 32'hCC800001); // -67108869
      convertSigned(64'h000000000400000B, 32'h4C800001); // 67108875
      convertSigned(64'hFFFFFFFFFBFFFFF5, 32'hCC800001); // -67108875
      convertSigned(64'h000000000400000C, 32'h4C800002); // 67108876
      convertSigned(64'hFFFFFFFFFBFFFFF4, 32'hCC800002); // -67108876
      convertSigned(64'h000000000400000D, 32'h4C800002); // 67108877
      convertSigned(64'hFFFFFFFFFBFFFFF3, 32'hCC800002); // -67108877
      convertSigned(64'h0000000008000007, 32'h4D000000); // 134217735
      convertSigned(64'hFFFFFFFFF7FFFFF9, 32'hCD000000); // -134217735
      convertSigned(64'h0000000008000008, 32'h4D000000); // 134217736
      convertSigned(64'hFFFFFFFFF7FFFFF8, 32'hCD000000); // -134217736
      convertSigned(64'h0000000008000009, 32'h4D000001); // 134217737
      convertSigned(64'hFFFFFFFFF7FFFFF7, 32'hCD000001); // -134217737
      convertSigned(64'h0000000008000017, 32'h4D000001); // 134217751
      convertSigned(64'hFFFFFFFFF7FFFFE9, 32'hCD000001); // -134217751
      convertSigned(64'h0000000008000018, 32'h4D000002); // 134217752
      convertSigned(64'hFFFFFFFFF7FFFFE8, 32'hCD000002); // -134217752
      convertSigned(64'h0000000008000019, 32'h4D000002); // 134217753
      convertSigned(64'hFFFFFFFFF7FFFFE7, 32'hCD000002); // -134217753
      convertSigned(64'h000000001000000F, 32'h4D800000); // 268435471
      convertSigned(64'hFFFFFFFFEFFFFFF1, 32'hCD800000); // -268435471
      convertSigned(64'h0000000010000010, 32'h4D800000); // 268435472
      convertSigned(64'hFFFFFFFFEFFFFFF0, 32'hCD800000); // -268435472
      convertSigned(64'h0000000010000011, 32'h4D800001); // 268435473
      convertSigned(64'hFFFFFFFFEFFFFFEF, 32'hCD800001); // -268435473
      convertSigned(64'h000000001000002F, 32'h4D800001); // 268435503
      convertSigned(64'hFFFFFFFFEFFFFFD1, 32'hCD800001); // -268435503
      convertSigned(64'h0000000010000030, 32'h4D800002); // 268435504
      convertSigned(64'hFFFFFFFFEFFFFFD0, 32'hCD800002); // -268435504
      convertSigned(64'h0000000010000031, 32'h4D800002); // 268435505
      convertSigned(64'hFFFFFFFFEFFFFFCF, 32'hCD800002); // -268435505
      convertSigned(64'h000000002000001F, 32'h4E000000); // 536870943
      convertSigned(64'hFFFFFFFFDFFFFFE1, 32'hCE000000); // -536870943
      convertSigned(64'h0000000020000020, 32'h4E000000); // 536870944
      convertSigned(64'hFFFFFFFFDFFFFFE0, 32'hCE000000); // -536870944
      convertSigned(64'h0000000020000021, 32'h4E000001); // 536870945
      convertSigned(64'hFFFFFFFFDFFFFFDF, 32'hCE000001); // -536870945
      convertSigned(64'h000000002000005F, 32'h4E000001); // 536871007
      convertSigned(64'hFFFFFFFFDFFFFFA1, 32'hCE000001); // -536871007
      convertSigned(64'h0000000020000060, 32'h4E000002); // 536871008
      convertSigned(64'hFFFFFFFFDFFFFFA0, 32'hCE000002); // -536871008
      convertSigned(64'h0000000020000061, 32'h4E000002); // 536871009
      convertSigned(64'hFFFFFFFFDFFFFF9F, 32'hCE000002); // -536871009
      convertSigned(64'h000000004000003F, 32'h4E800000); // 1073741887
      convertSigned(64'hFFFFFFFFBFFFFFC1, 32'hCE800000); // -1073741887
      convertSigned(64'h0000000040000040, 32'h4E800000); // 1073741888
      convertSigned(64'hFFFFFFFFBFFFFFC0, 32'hCE800000); // -1073741888
      convertSigned(64'h0000000040000041, 32'h4E800001); // 1073741889
      convertSigned(64'hFFFFFFFFBFFFFFBF, 32'hCE800001); // -1073741889
      convertSigned(64'h00000000400000BF, 32'h4E800001); // 1073742015
      convertSigned(64'hFFFFFFFFBFFFFF41, 32'hCE800001); // -1073742015
      convertSigned(64'h00000000400000C0, 32'h4E800002); // 1073742016
      convertSigned(64'hFFFFFFFFBFFFFF40, 32'hCE800002); // -1073742016
      convertSigned(64'h00000000400000C1, 32'h4E800002); // 1073742017
      convertSigned(64'hFFFFFFFFBFFFFF3F, 32'hCE800002); // -1073742017
      convertSigned(64'h000000008000007F, 32'h4F000000); // 2147483775
      convertSigned(64'hFFFFFFFF7FFFFF81, 32'hCF000000); // -2147483775
      convertSigned(64'h0000000080000080, 32'h4F000000); // 2147483776
      convertSigned(64'hFFFFFFFF7FFFFF80, 32'hCF000000); // -2147483776
      convertSigned(64'h0000000080000081, 32'h4F000001); // 2147483777
      convertSigned(64'hFFFFFFFF7FFFFF7F, 32'hCF000001); // -2147483777
      convertSigned(64'h000000008000017F, 32'h4F000001); // 2147484031
      convertSigned(64'hFFFFFFFF7FFFFE81, 32'hCF000001); // -2147484031
      convertSigned(64'h0000000080000180, 32'h4F000002); // 2147484032
      convertSigned(64'hFFFFFFFF7FFFFE80, 32'hCF000002); // -2147484032
      convertSigned(64'h0000000080000181, 32'h4F000002); // 2147484033
      convertSigned(64'hFFFFFFFF7FFFFE7F, 32'hCF000002); // -2147484033
      convertSigned(64'h00000001000000FF, 32'h4F800000); // 4294967551
      convertSigned(64'hFFFFFFFEFFFFFF01, 32'hCF800000); // -4294967551
      convertSigned(64'h0000000100000100, 32'h4F800000); // 4294967552
      convertSigned(64'hFFFFFFFEFFFFFF00, 32'hCF800000); // -4294967552
      convertSigned(64'h0000000100000101, 32'h4F800001); // 4294967553
      convertSigned(64'hFFFFFFFEFFFFFEFF, 32'hCF800001); // -4294967553
      convertSigned(64'h00000001000002FF, 32'h4F800001); // 4294968063
      convertSigned(64'hFFFFFFFEFFFFFD01, 32'hCF800001); // -4294968063
      convertSigned(64'h0000000100000300, 32'h4F800002); // 4294968064
      convertSigned(64'hFFFFFFFEFFFFFD00, 32'hCF800002); // -4294968064
      convertSigned(64'h0000000100000301, 32'h4F800002); // 4294968065
      convertSigned(64'hFFFFFFFEFFFFFCFF, 32'hCF800002); // -4294968065
      convertSigned(64'h00000002000001FF, 32'h50000000); // 8589935103
      convertSigned(64'hFFFFFFFDFFFFFE01, 32'hD0000000); // -8589935103
      convertSigned(64'h0000000200000200, 32'h50000000); // 8589935104
      convertSigned(64'hFFFFFFFDFFFFFE00, 32'hD0000000); // -8589935104
      convertSigned(64'h0000000200000201, 32'h50000001); // 8589935105
      convertSigned(64'hFFFFFFFDFFFFFDFF, 32'hD0000001); // -8589935105
      convertSigned(64'h00000002000005FF, 32'h50000001); // 8589936127
      convertSigned(64'hFFFFFFFDFFFFFA01, 32'hD0000001); // -8589936127
      convertSigned(64'h0000000200000600, 32'h50000002); // 8589936128
      convertSigned(64'hFFFFFFFDFFFFFA00, 32'hD0000002); // -8589936128
      convertSigned(64'h0000000200000601, 32'h50000002); // 8589936129
      convertSigned(64'hFFFFFFFDFFFFF9FF, 32'hD0000002); // -8589936129
      convertSigned(64'h00000004000003FF, 32'h50800000); // 17179870207
      convertSigned(64'hFFFFFFFBFFFFFC01, 32'hD0800000); // -17179870207
      convertSigned(64'h0000000400000400, 32'h50800000); // 17179870208
      convertSigned(64'hFFFFFFFBFFFFFC00, 32'hD0800000); // -17179870208
      convertSigned(64'h0000000400000401, 32'h50800001); // 17179870209
      convertSigned(64'hFFFFFFFBFFFFFBFF, 32'hD0800001); // -17179870209
      convertSigned(64'h0000000400000BFF, 32'h50800001); // 17179872255
      convertSigned(64'hFFFFFFFBFFFFF401, 32'hD0800001); // -17179872255
      convertSigned(64'h0000000400000C00, 32'h50800002); // 17179872256
      convertSigned(64'hFFFFFFFBFFFFF400, 32'hD0800002); // -17179872256
      convertSigned(64'h0000000400000C01, 32'h50800002); // 17179872257
      convertSigned(64'hFFFFFFFBFFFFF3FF, 32'hD0800002); // -17179872257
      convertSigned(64'h00000008000007FF, 32'h51000000); // 34359740415
      convertSigned(64'hFFFFFFF7FFFFF801, 32'hD1000000); // -34359740415
      convertSigned(64'h0000000800000800, 32'h51000000); // 34359740416
      convertSigned(64'hFFFFFFF7FFFFF800, 32'hD1000000); // -34359740416
      convertSigned(64'h0000000800000801, 32'h51000001); // 34359740417
      convertSigned(64'hFFFFFFF7FFFFF7FF, 32'hD1000001); // -34359740417
      convertSigned(64'h00000008000017FF, 32'h51000001); // 34359744511
      convertSigned(64'hFFFFFFF7FFFFE801, 32'hD1000001); // -34359744511
      convertSigned(64'h0000000800001800, 32'h51000002); // 34359744512
      convertSigned(64'hFFFFFFF7FFFFE800, 32'hD1000002); // -34359744512
      convertSigned(64'h0000000800001801, 32'h51000002); // 34359744513
      convertSigned(64'hFFFFFFF7FFFFE7FF, 32'hD1000002); // -34359744513
      convertSigned(64'h0000001000000FFF, 32'h51800000); // 68719480831
      convertSigned(64'hFFFFFFEFFFFFF001, 32'hD1800000); // -68719480831
      convertSigned(64'h0000001000001000, 32'h51800000); // 68719480832
      convertSigned(64'hFFFFFFEFFFFFF000, 32'hD1800000); // -68719480832
      convertSigned(64'h0000001000001001, 32'h51800001); // 68719480833
      convertSigned(64'hFFFFFFEFFFFFEFFF, 32'hD1800001); // -68719480833
      convertSigned(64'h0000001000002FFF, 32'h51800001); // 68719489023
      convertSigned(64'hFFFFFFEFFFFFD001, 32'hD1800001); // -68719489023
      convertSigned(64'h0000001000003000, 32'h51800002); // 68719489024
      convertSigned(64'hFFFFFFEFFFFFD000, 32'hD1800002); // -68719489024
      convertSigned(64'h0000001000003001, 32'h51800002); // 68719489025
      convertSigned(64'hFFFFFFEFFFFFCFFF, 32'hD1800002); // -68719489025
      convertSigned(64'h0000002000001FFF, 32'h52000000); // 137438961663
      convertSigned(64'hFFFFFFDFFFFFE001, 32'hD2000000); // -137438961663
      convertSigned(64'h0000002000002000, 32'h52000000); // 137438961664
      convertSigned(64'hFFFFFFDFFFFFE000, 32'hD2000000); // -137438961664
      convertSigned(64'h0000002000002001, 32'h52000001); // 137438961665
      convertSigned(64'hFFFFFFDFFFFFDFFF, 32'hD2000001); // -137438961665
      convertSigned(64'h0000002000005FFF, 32'h52000001); // 137438978047
      convertSigned(64'hFFFFFFDFFFFFA001, 32'hD2000001); // -137438978047
      convertSigned(64'h0000002000006000, 32'h52000002); // 137438978048
      convertSigned(64'hFFFFFFDFFFFFA000, 32'hD2000002); // -137438978048
      convertSigned(64'h0000002000006001, 32'h52000002); // 137438978049
      convertSigned(64'hFFFFFFDFFFFF9FFF, 32'hD2000002); // -137438978049
      convertSigned(64'h0000004000003FFF, 32'h52800000); // 274877923327
      convertSigned(64'hFFFFFFBFFFFFC001, 32'hD2800000); // -274877923327
      convertSigned(64'h0000004000004000, 32'h52800000); // 274877923328
      convertSigned(64'hFFFFFFBFFFFFC000, 32'hD2800000); // -274877923328
      convertSigned(64'h0000004000004001, 32'h52800001); // 274877923329
      convertSigned(64'hFFFFFFBFFFFFBFFF, 32'hD2800001); // -274877923329
      convertSigned(64'h000000400000BFFF, 32'h52800001); // 274877956095
      convertSigned(64'hFFFFFFBFFFFF4001, 32'hD2800001); // -274877956095
      convertSigned(64'h000000400000C000, 32'h52800002); // 274877956096
      convertSigned(64'hFFFFFFBFFFFF4000, 32'hD2800002); // -274877956096
      convertSigned(64'h000000400000C001, 32'h52800002); // 274877956097
      convertSigned(64'hFFFFFFBFFFFF3FFF, 32'hD2800002); // -274877956097
      convertSigned(64'h0000008000007FFF, 32'h53000000); // 549755846655
      convertSigned(64'hFFFFFF7FFFFF8001, 32'hD3000000); // -549755846655
      convertSigned(64'h0000008000008000, 32'h53000000); // 549755846656
      convertSigned(64'hFFFFFF7FFFFF8000, 32'hD3000000); // -549755846656
      convertSigned(64'h0000008000008001, 32'h53000001); // 549755846657
      convertSigned(64'hFFFFFF7FFFFF7FFF, 32'hD3000001); // -549755846657
      convertSigned(64'h0000008000017FFF, 32'h53000001); // 549755912191
      convertSigned(64'hFFFFFF7FFFFE8001, 32'hD3000001); // -549755912191
      convertSigned(64'h0000008000018000, 32'h53000002); // 549755912192
      convertSigned(64'hFFFFFF7FFFFE8000, 32'hD3000002); // -549755912192
      convertSigned(64'h0000008000018001, 32'h53000002); // 549755912193
      convertSigned(64'hFFFFFF7FFFFE7FFF, 32'hD3000002); // -549755912193
      convertSigned(64'h000001000000FFFF, 32'h53800000); // 1099511693311
      convertSigned(64'hFFFFFEFFFFFF0001, 32'hD3800000); // -1099511693311
      convertSigned(64'h0000010000010000, 32'h53800000); // 1099511693312
      convertSigned(64'hFFFFFEFFFFFF0000, 32'hD3800000); // -1099511693312
      convertSigned(64'h0000010000010001, 32'h53800001); // 1099511693313
      convertSigned(64'hFFFFFEFFFFFEFFFF, 32'hD3800001); // -1099511693313
      convertSigned(64'h000001000002FFFF, 32'h53800001); // 1099511824383
      convertSigned(64'hFFFFFEFFFFFD0001, 32'hD3800001); // -1099511824383
      convertSigned(64'h0000010000030000, 32'h53800002); // 1099511824384
      convertSigned(64'hFFFFFEFFFFFD0000, 32'hD3800002); // -1099511824384
      convertSigned(64'h0000010000030001, 32'h53800002); // 1099511824385
      convertSigned(64'hFFFFFEFFFFFCFFFF, 32'hD3800002); // -1099511824385
      convertSigned(64'h000002000001FFFF, 32'h54000000); // 2199023386623
      convertSigned(64'hFFFFFDFFFFFE0001, 32'hD4000000); // -2199023386623
      convertSigned(64'h0000020000020000, 32'h54000000); // 2199023386624
      convertSigned(64'hFFFFFDFFFFFE0000, 32'hD4000000); // -2199023386624
      convertSigned(64'h0000020000020001, 32'h54000001); // 2199023386625
      convertSigned(64'hFFFFFDFFFFFDFFFF, 32'hD4000001); // -2199023386625
      convertSigned(64'h000002000005FFFF, 32'h54000001); // 2199023648767
      convertSigned(64'hFFFFFDFFFFFA0001, 32'hD4000001); // -2199023648767
      convertSigned(64'h0000020000060000, 32'h54000002); // 2199023648768
      convertSigned(64'hFFFFFDFFFFFA0000, 32'hD4000002); // -2199023648768
      convertSigned(64'h0000020000060001, 32'h54000002); // 2199023648769
      convertSigned(64'hFFFFFDFFFFF9FFFF, 32'hD4000002); // -2199023648769
      convertSigned(64'h000004000003FFFF, 32'h54800000); // 4398046773247
      convertSigned(64'hFFFFFBFFFFFC0001, 32'hD4800000); // -4398046773247
      convertSigned(64'h0000040000040000, 32'h54800000); // 4398046773248
      convertSigned(64'hFFFFFBFFFFFC0000, 32'hD4800000); // -4398046773248
      convertSigned(64'h0000040000040001, 32'h54800001); // 4398046773249
      convertSigned(64'hFFFFFBFFFFFBFFFF, 32'hD4800001); // -4398046773249
      convertSigned(64'h00000400000BFFFF, 32'h54800001); // 4398047297535
      convertSigned(64'hFFFFFBFFFFF40001, 32'hD4800001); // -4398047297535
      convertSigned(64'h00000400000C0000, 32'h54800002); // 4398047297536
      convertSigned(64'hFFFFFBFFFFF40000, 32'hD4800002); // -4398047297536
      convertSigned(64'h00000400000C0001, 32'h54800002); // 4398047297537
      convertSigned(64'hFFFFFBFFFFF3FFFF, 32'hD4800002); // -4398047297537
      convertSigned(64'h000008000007FFFF, 32'h55000000); // 8796093546495
      convertSigned(64'hFFFFF7FFFFF80001, 32'hD5000000); // -8796093546495
      convertSigned(64'h0000080000080000, 32'h55000000); // 8796093546496
      convertSigned(64'hFFFFF7FFFFF80000, 32'hD5000000); // -8796093546496
      convertSigned(64'h0000080000080001, 32'h55000001); // 8796093546497
      convertSigned(64'hFFFFF7FFFFF7FFFF, 32'hD5000001); // -8796093546497
      convertSigned(64'h000008000017FFFF, 32'h55000001); // 8796094595071
      convertSigned(64'hFFFFF7FFFFE80001, 32'hD5000001); // -8796094595071
      convertSigned(64'h0000080000180000, 32'h55000002); // 8796094595072
      convertSigned(64'hFFFFF7FFFFE80000, 32'hD5000002); // -8796094595072
      convertSigned(64'h0000080000180001, 32'h55000002); // 8796094595073
      convertSigned(64'hFFFFF7FFFFE7FFFF, 32'hD5000002); // -8796094595073
      convertSigned(64'h00001000000FFFFF, 32'h55800000); // 17592187092991
      convertSigned(64'hFFFFEFFFFFF00001, 32'hD5800000); // -17592187092991
      convertSigned(64'h0000100000100000, 32'h55800000); // 17592187092992
      convertSigned(64'hFFFFEFFFFFF00000, 32'hD5800000); // -17592187092992
      convertSigned(64'h0000100000100001, 32'h55800001); // 17592187092993
      convertSigned(64'hFFFFEFFFFFEFFFFF, 32'hD5800001); // -17592187092993
      convertSigned(64'h00001000002FFFFF, 32'h55800001); // 17592189190143
      convertSigned(64'hFFFFEFFFFFD00001, 32'hD5800001); // -17592189190143
      convertSigned(64'h0000100000300000, 32'h55800002); // 17592189190144
      convertSigned(64'hFFFFEFFFFFD00000, 32'hD5800002); // -17592189190144
      convertSigned(64'h0000100000300001, 32'h55800002); // 17592189190145
      convertSigned(64'hFFFFEFFFFFCFFFFF, 32'hD5800002); // -17592189190145
      convertSigned(64'h00002000001FFFFF, 32'h56000000); // 35184374185983
      convertSigned(64'hFFFFDFFFFFE00001, 32'hD6000000); // -35184374185983
      convertSigned(64'h0000200000200000, 32'h56000000); // 35184374185984
      convertSigned(64'hFFFFDFFFFFE00000, 32'hD6000000); // -35184374185984
      convertSigned(64'h0000200000200001, 32'h56000001); // 35184374185985
      convertSigned(64'hFFFFDFFFFFDFFFFF, 32'hD6000001); // -35184374185985
      convertSigned(64'h00002000005FFFFF, 32'h56000001); // 35184378380287
      convertSigned(64'hFFFFDFFFFFA00001, 32'hD6000001); // -35184378380287
      convertSigned(64'h0000200000600000, 32'h56000002); // 35184378380288
      convertSigned(64'hFFFFDFFFFFA00000, 32'hD6000002); // -35184378380288
      convertSigned(64'h0000200000600001, 32'h56000002); // 35184378380289
      convertSigned(64'hFFFFDFFFFF9FFFFF, 32'hD6000002); // -35184378380289
      convertSigned(64'h00004000003FFFFF, 32'h56800000); // 70368748371967
      convertSigned(64'hFFFFBFFFFFC00001, 32'hD6800000); // -70368748371967
      convertSigned(64'h0000400000400000, 32'h56800000); // 70368748371968
      convertSigned(64'hFFFFBFFFFFC00000, 32'hD6800000); // -70368748371968
      convertSigned(64'h0000400000400001, 32'h56800001); // 70368748371969
      convertSigned(64'hFFFFBFFFFFBFFFFF, 32'hD6800001); // -70368748371969
      convertSigned(64'h0000400000BFFFFF, 32'h56800001); // 70368756760575
      convertSigned(64'hFFFFBFFFFF400001, 32'hD6800001); // -70368756760575
      convertSigned(64'h0000400000C00000, 32'h56800002); // 70368756760576
      convertSigned(64'hFFFFBFFFFF400000, 32'hD6800002); // -70368756760576
      convertSigned(64'h0000400000C00001, 32'h56800002); // 70368756760577
      convertSigned(64'hFFFFBFFFFF3FFFFF, 32'hD6800002); // -70368756760577
      convertSigned(64'h00008000007FFFFF, 32'h57000000); // 140737496743935
      convertSigned(64'hFFFF7FFFFF800001, 32'hD7000000); // -140737496743935
      convertSigned(64'h0000800000800000, 32'h57000000); // 140737496743936
      convertSigned(64'hFFFF7FFFFF800000, 32'hD7000000); // -140737496743936
      convertSigned(64'h0000800000800001, 32'h57000001); // 140737496743937
      convertSigned(64'hFFFF7FFFFF7FFFFF, 32'hD7000001); // -140737496743937
      convertSigned(64'h00008000017FFFFF, 32'h57000001); // 140737513521151
      convertSigned(64'hFFFF7FFFFE800001, 32'hD7000001); // -140737513521151
      convertSigned(64'h0000800001800000, 32'h57000002); // 140737513521152
      convertSigned(64'hFFFF7FFFFE800000, 32'hD7000002); // -140737513521152
      convertSigned(64'h0000800001800001, 32'h57000002); // 140737513521153
      convertSigned(64'hFFFF7FFFFE7FFFFF, 32'hD7000002); // -140737513521153
      convertSigned(64'h0001000000FFFFFF, 32'h57800000); // 281474993487871
      convertSigned(64'hFFFEFFFFFF000001, 32'hD7800000); // -281474993487871
      convertSigned(64'h0001000001000000, 32'h57800000); // 281474993487872
      convertSigned(64'hFFFEFFFFFF000000, 32'hD7800000); // -281474993487872
      convertSigned(64'h0001000001000001, 32'h57800001); // 281474993487873
      convertSigned(64'hFFFEFFFFFEFFFFFF, 32'hD7800001); // -281474993487873
      convertSigned(64'h0001000002FFFFFF, 32'h57800001); // 281475027042303
      convertSigned(64'hFFFEFFFFFD000001, 32'hD7800001); // -281475027042303
      convertSigned(64'h0001000003000000, 32'h57800002); // 281475027042304
      convertSigned(64'hFFFEFFFFFD000000, 32'hD7800002); // -281475027042304
      convertSigned(64'h0001000003000001, 32'h57800002); // 281475027042305
      convertSigned(64'hFFFEFFFFFCFFFFFF, 32'hD7800002); // -281475027042305
      convertSigned(64'h0002000001FFFFFF, 32'h58000000); // 562949986975743
      convertSigned(64'hFFFDFFFFFE000001, 32'hD8000000); // -562949986975743
      convertSigned(64'h0002000002000000, 32'h58000000); // 562949986975744
      convertSigned(64'hFFFDFFFFFE000000, 32'hD8000000); // -562949986975744
      convertSigned(64'h0002000002000001, 32'h58000001); // 562949986975745
      convertSigned(64'hFFFDFFFFFDFFFFFF, 32'hD8000001); // -562949986975745
      convertSigned(64'h0002000005FFFFFF, 32'h58000001); // 562950054084607
      convertSigned(64'hFFFDFFFFFA000001, 32'hD8000001); // -562950054084607
      convertSigned(64'h0002000006000000, 32'h58000002); // 562950054084608
      convertSigned(64'hFFFDFFFFFA000000, 32'hD8000002); // -562950054084608
      convertSigned(64'h0002000006000001, 32'h58000002); // 562950054084609
      convertSigned(64'hFFFDFFFFF9FFFFFF, 32'hD8000002); // -562950054084609
      convertSigned(64'h0004000003FFFFFF, 32'h58800000); // 1125899973951487
      convertSigned(64'hFFFBFFFFFC000001, 32'hD8800000); // -1125899973951487
      convertSigned(64'h0004000004000000, 32'h58800000); // 1125899973951488
      convertSigned(64'hFFFBFFFFFC000000, 32'hD8800000); // -1125899973951488
      convertSigned(64'h0004000004000001, 32'h58800001); // 1125899973951489
      convertSigned(64'hFFFBFFFFFBFFFFFF, 32'hD8800001); // -1125899973951489
      convertSigned(64'h000400000BFFFFFF, 32'h58800001); // 1125900108169215
      convertSigned(64'hFFFBFFFFF4000001, 32'hD8800001); // -1125900108169215
      convertSigned(64'h000400000C000000, 32'h58800002); // 1125900108169216
      convertSigned(64'hFFFBFFFFF4000000, 32'hD8800002); // -1125900108169216
      convertSigned(64'h000400000C000001, 32'h58800002); // 1125900108169217
      convertSigned(64'hFFFBFFFFF3FFFFFF, 32'hD8800002); // -1125900108169217
      convertSigned(64'h0008000007FFFFFF, 32'h59000000); // 2251799947902975
      convertSigned(64'hFFF7FFFFF8000001, 32'hD9000000); // -2251799947902975
      convertSigned(64'h0008000008000000, 32'h59000000); // 2251799947902976
      convertSigned(64'hFFF7FFFFF8000000, 32'hD9000000); // -2251799947902976
      convertSigned(64'h0008000008000001, 32'h59000001); // 2251799947902977
      convertSigned(64'hFFF7FFFFF7FFFFFF, 32'hD9000001); // -2251799947902977
      convertSigned(64'h0008000017FFFFFF, 32'h59000001); // 2251800216338431
      convertSigned(64'hFFF7FFFFE8000001, 32'hD9000001); // -2251800216338431
      convertSigned(64'h0008000018000000, 32'h59000002); // 2251800216338432
      convertSigned(64'hFFF7FFFFE8000000, 32'hD9000002); // -2251800216338432
      convertSigned(64'h0008000018000001, 32'h59000002); // 2251800216338433
      convertSigned(64'hFFF7FFFFE7FFFFFF, 32'hD9000002); // -2251800216338433
      convertSigned(64'h001000000FFFFFFF, 32'h59800000); // 4503599895805951
      convertSigned(64'hFFEFFFFFF0000001, 32'hD9800000); // -4503599895805951
      convertSigned(64'h0010000010000000, 32'h59800000); // 4503599895805952
      convertSigned(64'hFFEFFFFFF0000000, 32'hD9800000); // -4503599895805952
      convertSigned(64'h0010000010000001, 32'h59800001); // 4503599895805953
      convertSigned(64'hFFEFFFFFEFFFFFFF, 32'hD9800001); // -4503599895805953
      convertSigned(64'h001000002FFFFFFF, 32'h59800001); // 4503600432676863
      convertSigned(64'hFFEFFFFFD0000001, 32'hD9800001); // -4503600432676863
      convertSigned(64'h0010000030000000, 32'h59800002); // 4503600432676864
      convertSigned(64'hFFEFFFFFD0000000, 32'hD9800002); // -4503600432676864
      convertSigned(64'h0010000030000001, 32'h59800002); // 4503600432676865
      convertSigned(64'hFFEFFFFFCFFFFFFF, 32'hD9800002); // -4503600432676865
      convertSigned(64'h002000001FFFFFFF, 32'h5A000000); // 9007199791611903
      convertSigned(64'hFFDFFFFFE0000001, 32'hDA000000); // -9007199791611903
      convertSigned(64'h0020000020000000, 32'h5A000000); // 9007199791611904
      convertSigned(64'hFFDFFFFFE0000000, 32'hDA000000); // -9007199791611904
      convertSigned(64'h0020000020000001, 32'h5A000001); // 9007199791611905
      convertSigned(64'hFFDFFFFFDFFFFFFF, 32'hDA000001); // -9007199791611905
      convertSigned(64'h002000005FFFFFFF, 32'h5A000001); // 9007200865353727
      convertSigned(64'hFFDFFFFFA0000001, 32'hDA000001); // -9007200865353727
      convertSigned(64'h0020000060000000, 32'h5A000002); // 9007200865353728
      convertSigned(64'hFFDFFFFFA0000000, 32'hDA000002); // -9007200865353728
      convertSigned(64'h0020000060000001, 32'h5A000002); // 9007200865353729
      convertSigned(64'hFFDFFFFF9FFFFFFF, 32'hDA000002); // -9007200865353729
      convertSigned(64'h004000003FFFFFFF, 32'h5A800000); // 18014399583223807
      convertSigned(64'hFFBFFFFFC0000001, 32'hDA800000); // -18014399583223807
      convertSigned(64'h0040000040000000, 32'h5A800000); // 18014399583223808
      convertSigned(64'hFFBFFFFFC0000000, 32'hDA800000); // -18014399583223808
      convertSigned(64'h0040000040000001, 32'h5A800001); // 18014399583223809
      convertSigned(64'hFFBFFFFFBFFFFFFF, 32'hDA800001); // -18014399583223809
      convertSigned(64'h00400000BFFFFFFF, 32'h5A800001); // 18014401730707455
      convertSigned(64'hFFBFFFFF40000001, 32'hDA800001); // -18014401730707455
      convertSigned(64'h00400000C0000000, 32'h5A800002); // 18014401730707456
      convertSigned(64'hFFBFFFFF40000000, 32'hDA800002); // -18014401730707456
      convertSigned(64'h00400000C0000001, 32'h5A800002); // 18014401730707457
      convertSigned(64'hFFBFFFFF3FFFFFFF, 32'hDA800002); // -18014401730707457
      convertSigned(64'h008000007FFFFFFF, 32'h5B000000); // 36028799166447615
      convertSigned(64'hFF7FFFFF80000001, 32'hDB000000); // -36028799166447615
      convertSigned(64'h0080000080000000, 32'h5B000000); // 36028799166447616
      convertSigned(64'hFF7FFFFF80000000, 32'hDB000000); // -36028799166447616
      convertSigned(64'h0080000080000001, 32'h5B000001); // 36028799166447617
      convertSigned(64'hFF7FFFFF7FFFFFFF, 32'hDB000001); // -36028799166447617
      convertSigned(64'h008000017FFFFFFF, 32'h5B000001); // 36028803461414911
      convertSigned(64'hFF7FFFFE80000001, 32'hDB000001); // -36028803461414911
      convertSigned(64'h0080000180000000, 32'h5B000002); // 36028803461414912
      convertSigned(64'hFF7FFFFE80000000, 32'hDB000002); // -36028803461414912
      convertSigned(64'h0080000180000001, 32'h5B000002); // 36028803461414913
      convertSigned(64'hFF7FFFFE7FFFFFFF, 32'hDB000002); // -36028803461414913
      convertSigned(64'h01000000FFFFFFFF, 32'h5B800000); // 72057598332895231
      convertSigned(64'hFEFFFFFF00000001, 32'hDB800000); // -72057598332895231
      convertSigned(64'h0100000100000000, 32'h5B800000); // 72057598332895232
      convertSigned(64'hFEFFFFFF00000000, 32'hDB800000); // -72057598332895232
      convertSigned(64'h0100000100000001, 32'h5B800001); // 72057598332895233
      convertSigned(64'hFEFFFFFEFFFFFFFF, 32'hDB800001); // -72057598332895233
      convertSigned(64'h01000002FFFFFFFF, 32'h5B800001); // 72057606922829823
      convertSigned(64'hFEFFFFFD00000001, 32'hDB800001); // -72057606922829823
      convertSigned(64'h0100000300000000, 32'h5B800002); // 72057606922829824
      convertSigned(64'hFEFFFFFD00000000, 32'hDB800002); // -72057606922829824
      convertSigned(64'h0100000300000001, 32'h5B800002); // 72057606922829825
      convertSigned(64'hFEFFFFFCFFFFFFFF, 32'hDB800002); // -72057606922829825
      convertSigned(64'h02000001FFFFFFFF, 32'h5C000000); // 144115196665790463
      convertSigned(64'hFDFFFFFE00000001, 32'hDC000000); // -144115196665790463
      convertSigned(64'h0200000200000000, 32'h5C000000); // 144115196665790464
      convertSigned(64'hFDFFFFFE00000000, 32'hDC000000); // -144115196665790464
      convertSigned(64'h0200000200000001, 32'h5C000001); // 144115196665790465
      convertSigned(64'hFDFFFFFDFFFFFFFF, 32'hDC000001); // -144115196665790465
      convertSigned(64'h02000005FFFFFFFF, 32'h5C000001); // 144115213845659647
      convertSigned(64'hFDFFFFFA00000001, 32'hDC000001); // -144115213845659647
      convertSigned(64'h0200000600000000, 32'h5C000002); // 144115213845659648
      convertSigned(64'hFDFFFFFA00000000, 32'hDC000002); // -144115213845659648
      convertSigned(64'h0200000600000001, 32'h5C000002); // 144115213845659649
      convertSigned(64'hFDFFFFF9FFFFFFFF, 32'hDC000002); // -144115213845659649
      convertSigned(64'h04000003FFFFFFFF, 32'h5C800000); // 288230393331580927
      convertSigned(64'hFBFFFFFC00000001, 32'hDC800000); // -288230393331580927
      convertSigned(64'h0400000400000000, 32'h5C800000); // 288230393331580928
      convertSigned(64'hFBFFFFFC00000000, 32'hDC800000); // -288230393331580928
      convertSigned(64'h0400000400000001, 32'h5C800001); // 288230393331580929
      convertSigned(64'hFBFFFFFBFFFFFFFF, 32'hDC800001); // -288230393331580929
      convertSigned(64'h0400000BFFFFFFFF, 32'h5C800001); // 288230427691319295
      convertSigned(64'hFBFFFFF400000001, 32'hDC800001); // -288230427691319295
      convertSigned(64'h0400000C00000000, 32'h5C800002); // 288230427691319296
      convertSigned(64'hFBFFFFF400000000, 32'hDC800002); // -288230427691319296
      convertSigned(64'h0400000C00000001, 32'h5C800002); // 288230427691319297
      convertSigned(64'hFBFFFFF3FFFFFFFF, 32'hDC800002); // -288230427691319297
      convertSigned(64'h08000007FFFFFFFF, 32'h5D000000); // 576460786663161855
      convertSigned(64'hF7FFFFF800000001, 32'hDD000000); // -576460786663161855
      convertSigned(64'h0800000800000000, 32'h5D000000); // 576460786663161856
      convertSigned(64'hF7FFFFF800000000, 32'hDD000000); // -576460786663161856
      convertSigned(64'h0800000800000001, 32'h5D000001); // 576460786663161857
      convertSigned(64'hF7FFFFF7FFFFFFFF, 32'hDD000001); // -576460786663161857
      convertSigned(64'h08000017FFFFFFFF, 32'h5D000001); // 576460855382638591
      convertSigned(64'hF7FFFFE800000001, 32'hDD000001); // -576460855382638591
      convertSigned(64'h0800001800000000, 32'h5D000002); // 576460855382638592
      convertSigned(64'hF7FFFFE800000000, 32'hDD000002); // -576460855382638592
      convertSigned(64'h0800001800000001, 32'h5D000002); // 576460855382638593
      convertSigned(64'hF7FFFFE7FFFFFFFF, 32'hDD000002); // -576460855382638593
      convertSigned(64'h1000000FFFFFFFFF, 32'h5D800000); // 1152921573326323711
      convertSigned(64'hEFFFFFF000000001, 32'hDD800000); // -1152921573326323711
      convertSigned(64'h1000001000000000, 32'h5D800000); // 1152921573326323712
      convertSigned(64'hEFFFFFF000000000, 32'hDD800000); // -1152921573326323712
      convertSigned(64'h1000001000000001, 32'h5D800001); // 1152921573326323713
      convertSigned(64'hEFFFFFEFFFFFFFFF, 32'hDD800001); // -1152921573326323713
      convertSigned(64'h1000002FFFFFFFFF, 32'h5D800001); // 1152921710765277183
      convertSigned(64'hEFFFFFD000000001, 32'hDD800001); // -1152921710765277183
      convertSigned(64'h1000003000000000, 32'h5D800002); // 1152921710765277184
      convertSigned(64'hEFFFFFD000000000, 32'hDD800002); // -1152921710765277184
      convertSigned(64'h1000003000000001, 32'h5D800002); // 1152921710765277185
      convertSigned(64'hEFFFFFCFFFFFFFFF, 32'hDD800002); // -1152921710765277185
      convertSigned(64'h2000001FFFFFFFFF, 32'h5E000000); // 2305843146652647423
      convertSigned(64'hDFFFFFE000000001, 32'hDE000000); // -2305843146652647423
      convertSigned(64'h2000002000000000, 32'h5E000000); // 2305843146652647424
      convertSigned(64'hDFFFFFE000000000, 32'hDE000000); // -2305843146652647424
      convertSigned(64'h2000002000000001, 32'h5E000001); // 2305843146652647425
      convertSigned(64'hDFFFFFDFFFFFFFFF, 32'hDE000001); // -2305843146652647425
      convertSigned(64'h2000005FFFFFFFFF, 32'h5E000001); // 2305843421530554367
      convertSigned(64'hDFFFFFA000000001, 32'hDE000001); // -2305843421530554367
      convertSigned(64'h2000006000000000, 32'h5E000002); // 2305843421530554368
      convertSigned(64'hDFFFFFA000000000, 32'hDE000002); // -2305843421530554368
      convertSigned(64'h2000006000000001, 32'h5E000002); // 2305843421530554369
      convertSigned(64'hDFFFFF9FFFFFFFFF, 32'hDE000002); // -2305843421530554369
      convertSigned(64'h4000003FFFFFFFFF, 32'h5E800000); // 4611686293305294847
      convertSigned(64'hBFFFFFC000000001, 32'hDE800000); // -4611686293305294847
      convertSigned(64'h4000004000000000, 32'h5E800000); // 4611686293305294848
      convertSigned(64'hBFFFFFC000000000, 32'hDE800000); // -4611686293305294848
      convertSigned(64'h4000004000000001, 32'h5E800001); // 4611686293305294849
      convertSigned(64'hBFFFFFBFFFFFFFFF, 32'hDE800001); // -4611686293305294849
      convertSigned(64'h400000BFFFFFFFFF, 32'h5E800001); // 4611686843061108735
      convertSigned(64'hBFFFFF4000000001, 32'hDE800001); // -4611686843061108735
      convertSigned(64'h400000C000000000, 32'h5E800002); // 4611686843061108736
      convertSigned(64'hBFFFFF4000000000, 32'hDE800002); // -4611686843061108736
      convertSigned(64'h400000C000000001, 32'h5E800002); // 4611686843061108737
      convertSigned(64'hBFFFFF3FFFFFFFFF, 32'hDE800002); // -4611686843061108737
      
      // random signed test cases
      convertSigned(64'h8000000000000000, 32'hDF000000); // -9223372036854775808
      convertSigned(64'hFFFFFFFFFFC00000, 32'hCA800000); // -4194304
      convertSigned(64'hFFFFFFFFFF800000, 32'hCB000000); // -8388608
      convertSigned(64'hFFFFFFFFFF000000, 32'hCB800000); // -16777216
      convertSigned(64'hFFFFFFFFFF800000, 32'hCB000000); // -8388608
      convertSigned(64'hFFFFFFFFFF000000, 32'hCB800000); // -16777216
      convertSigned(64'hFFFFFFFFFE000000, 32'hCC000000); // -33554432
      convertSigned(64'hFFFFFFFFFFF0BDC0, 32'hC9742400); // -1000000
      convertSigned(64'hFFFFFFFFFFFFFFF6, 32'hC1200000); // -10
      convertSigned(64'hFFFFFFFFFFFFFFFF, 32'hBF800000); // -1
      convertSigned(64'h0000000000000000, 32'h00000000); // 0
      convertSigned(64'h0000000000000001, 32'h3F800000); // 1
      convertSigned(64'h000000000000000A, 32'h41200000); // 10
      convertSigned(64'h00000000000F4240, 32'h49742400); // 1000000
      convertSigned(64'h0000000000400000, 32'h4A800000); // 4194304
      convertSigned(64'h0000000000800000, 32'h4B000000); // 8388608
      convertSigned(64'h0000000001000000, 32'h4B800000); // 16777216
      convertSigned(64'h0000000000800000, 32'h4B000000); // 8388608
      convertSigned(64'h0000000001000000, 32'h4B800000); // 16777216
      convertSigned(64'h0000000002000000, 32'h4C000000); // 33554432
      convertSigned(64'h7FFFFFFFFFFFFFFF, 32'h5F000000); // 9223372036854775807
      convertSigned(64'h1649EC5F2C93D800, 32'h5DB24F63); // 1606074635648227328
      convertSigned(64'h00628499D2C50930, 32'h5AC50934); // 27730343918635312
      convertSigned(64'hFFFCA6DB8BBCE72D, 32'hD856491D); // -942438034381011
      convertSigned(64'h0000603A666CC074, 32'h56C074CD); // 105803942772852
      convertSigned(64'h00000B066DFFCDE8, 32'h553066E0); // 12122243190248
      convertSigned(64'h000012BCAF986F73, 32'h5595E57D); // 20601609154419
      convertSigned(64'hFFFFF5DE3522ECA2, 32'hD5221CAE); // -11140253684574
      convertSigned(64'h0000000E76D1A81C, 32'h51676D1B); // 62122993692
      convertSigned(64'h000000E9ACDA7B0B, 32'h5369ACDA); // 1003627379467
      convertSigned(64'h0000003C755A895B, 32'h5271D56A); // 259666905435
      convertSigned(64'hFFFFFF97EEA746C8, 32'hD2D022B1); // -446967626040
      convertSigned(64'h00000036548BF440, 32'h52595230); // 233346692160
      convertSigned(64'hFFFFFFFDEDAC61A7, 32'hD00494E8); // -8897404505
      convertSigned(64'hFFFFFFEDB1026F5A, 32'hD19277ED); // -78634651814
      convertSigned(64'h00000002DA25202E, 32'h50368948); // 12249800750
      convertSigned(64'hFFFFFFF8E9754F82, 32'hD0E2D156); // -30442958974
      convertSigned(64'hFFFFFFFDC08A7D41, 32'hD00FDD61); // -9654600383
      convertSigned(64'hFFFFFFFE2632103E, 32'hCFECE6F8); // -7949119426
      convertSigned(64'hFFFFFFFF2ED4D575, 32'hCF512B2B); // -3509267083
      convertSigned(64'h0000000016013B6C, 32'h4DB009DB); // 369179500
      convertSigned(64'hFFFFFFFFF36EDFDF, 32'hCD491202); // -210837537
      convertSigned(64'h000000003A7EF726, 32'h4E69FBDD); // 981399334
      convertSigned(64'h0000000030F3B575, 32'h4E43CED6); // 821278069
      convertSigned(64'hFFFFFFFFBC2D6179, 32'hCE87A53D); // -1137876615
      convertSigned(64'h00000000044A82BD, 32'h4C895058); // 71991997
      convertSigned(64'h000000001ED47D03, 32'h4DF6A3E8); // 517242115
      convertSigned(64'h000000002CBAE665, 32'h4E32EB9A); // 750446181
      convertSigned(64'hFFFFFFFFFE7E3C44, 32'hCBC0E1DE); // -25281468
      convertSigned(64'hFFFFFFFFFE199748, 32'hCBF3345C); // -31877304
      convertSigned(64'h000000000F092860, 32'h4D709286); // 252258400
      convertSigned(64'hFFFFFFFFF20369EF, 32'hCD5FC961); // -234657297
      convertSigned(64'h0000000004254347, 32'h4C84A869); // 69550919
      convertSigned(64'h0000000002506399, 32'h4C1418E6); // 38822809
      convertSigned(64'hFFFFFFFFF8F9BB42, 32'hCCE0C898); // -117851326
      convertSigned(64'hFFFFFFFFFF859A87, 32'hCAF4CAF2); // -8021369
      convertSigned(64'h00000000067A0D80, 32'h4CCF41B0); // 108662144
           
      convertSigned(64'h00000000067A0D80, 32'h4CCF41B0); // 108662144
      convertSigned(64'h00000000067A0D81, 32'h4CCF41B0); // 108662145
      convertSigned(64'h00000000067A0D82, 32'h4CCF41B0); // 108662146
      convertSigned(64'h00000000067A0D83, 32'h4CCF41B0); // 108662147
      convertSigned(64'h00000000067A0D84, 32'h4CCF41B0); // 108662148
      convertSigned(64'h00000000067A0D85, 32'h4CCF41B1); // 108662149
      convertSigned(64'h00000000067A0D86, 32'h4CCF41B1); // 108662150
      
      convertSigned(64'h000000000244D9BA, 32'h4C11366E); // 38066618
      convertSigned(64'hFFFFFFFFFDBB2646, 32'hCC11366E); // -38066618
      convertSigned(64'h00000000032DFBF4, 32'h4C4B7EFD); // 53345268
      convertSigned(64'hFFFFFFFFFC274CE5, 32'hCC762CC7); // -64533275
      convertSigned(64'hFFFFFFFFFEBCEB13, 32'hCBA18A76); // -21173485
      convertSigned(64'hFFFFFFFFFE63AE1D, 32'hCBCE28F2); // -27021795
      convertSigned(64'hFFFFFFFFFFBFE5D8, 32'hCA803450); // -4201000
      convertSigned(64'h000000000027F234, 32'h4A1FC8D0); // 2617908
      convertSigned(64'hFFFFFFFFFFC45AB0, 32'hCA6E9540); // -3908944
      convertSigned(64'hFFFFFFFFFF66D0D0, 32'hCB192F30); // -10039088
      convertSigned(64'hFFFFFFFFFF95030F, 32'hCAD5F9E2); // -7011569
      convertSigned(64'hFFFFFFFFFFD50864, 32'hCA2BDE70); // -2815900
      convertSigned(64'h0000000000AB9A8F, 32'h4B2B9A8F); // 11246223
      convertSigned(64'hFFFFFFFFFF99C83E, 32'hCACC6F84); // -6698946
      convertSigned(64'h00000000004B85AB, 32'h4A970B56); // 4949419
      
    end
    `uvm_info("LABEL", "Finished run phase.", UVM_HIGH);
    phase.drop_objection(this);
  endtask: run_phase
  
endclass

//-----------
// module top
//-----------
module top;

  bit clk;
  env environment;
  IntToFloat dut(.clk (clk));

  initial begin
    environment = new("env");
    // Put the interface into the resource database.
    uvm_resource_db#(virtual IntToFloat_IF)::set("env",
      "IntToFloat_IF", dut.IntToFloat_IF0);
    clk = 0;
    run_test();
  end
  
  initial begin
    forever begin
      #(50) clk = ~clk;
    end
  end
  
  initial begin
    // Dump waves
    $dumpvars(0, top);
  end
  
endmodule